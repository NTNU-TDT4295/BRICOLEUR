module FIFO( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input  [15:0] io_dataIn, // @[:@6.4]
  output [15:0] io_dataOut // @[:@6.4]
);
  reg [15:0] _T_11; // @[FIFO.scala 14:16:@8.4]
  reg [31:0] _RAND_0;
  assign io_dataOut = _T_11; // @[FIFO.scala 22:14:@9.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_11 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_11 <= 16'sh0;
    end else begin
      _T_11 <= io_dataIn;
    end
  end
endmodule
module FIFO_2( // @[:@21.2]
  input         clock, // @[:@22.4]
  input         reset, // @[:@23.4]
  input  [15:0] io_dataIn, // @[:@24.4]
  output [15:0] io_dataOut // @[:@24.4]
);
  reg [15:0] _T_11; // @[FIFO.scala 14:16:@26.4]
  reg [31:0] _RAND_0;
  reg [15:0] _T_14; // @[FIFO.scala 14:16:@27.4]
  reg [31:0] _RAND_1;
  reg [15:0] _T_17; // @[FIFO.scala 14:16:@28.4]
  reg [31:0] _RAND_2;
  reg [15:0] _T_20; // @[FIFO.scala 14:16:@29.4]
  reg [31:0] _RAND_3;
  reg [15:0] _T_23; // @[FIFO.scala 14:16:@30.4]
  reg [31:0] _RAND_4;
  reg [15:0] _T_26; // @[FIFO.scala 14:16:@31.4]
  reg [31:0] _RAND_5;
  reg [15:0] _T_29; // @[FIFO.scala 14:16:@32.4]
  reg [31:0] _RAND_6;
  reg [15:0] _T_32; // @[FIFO.scala 14:16:@33.4]
  reg [31:0] _RAND_7;
  reg [15:0] _T_35; // @[FIFO.scala 14:16:@34.4]
  reg [31:0] _RAND_8;
  reg [15:0] _T_38; // @[FIFO.scala 14:16:@35.4]
  reg [31:0] _RAND_9;
  reg [15:0] _T_41; // @[FIFO.scala 14:16:@36.4]
  reg [31:0] _RAND_10;
  reg [15:0] _T_44; // @[FIFO.scala 14:16:@37.4]
  reg [31:0] _RAND_11;
  reg [15:0] _T_47; // @[FIFO.scala 14:16:@38.4]
  reg [31:0] _RAND_12;
  reg [15:0] _T_50; // @[FIFO.scala 14:16:@39.4]
  reg [31:0] _RAND_13;
  reg [15:0] _T_53; // @[FIFO.scala 14:16:@40.4]
  reg [31:0] _RAND_14;
  reg [15:0] _T_56; // @[FIFO.scala 14:16:@41.4]
  reg [31:0] _RAND_15;
  reg [15:0] _T_59; // @[FIFO.scala 14:16:@42.4]
  reg [31:0] _RAND_16;
  reg [15:0] _T_62; // @[FIFO.scala 14:16:@43.4]
  reg [31:0] _RAND_17;
  reg [15:0] _T_65; // @[FIFO.scala 14:16:@44.4]
  reg [31:0] _RAND_18;
  reg [15:0] _T_68; // @[FIFO.scala 14:16:@45.4]
  reg [31:0] _RAND_19;
  reg [15:0] _T_71; // @[FIFO.scala 14:16:@46.4]
  reg [31:0] _RAND_20;
  reg [15:0] _T_74; // @[FIFO.scala 14:16:@47.4]
  reg [31:0] _RAND_21;
  reg [15:0] _T_77; // @[FIFO.scala 14:16:@48.4]
  reg [31:0] _RAND_22;
  reg [15:0] _T_80; // @[FIFO.scala 14:16:@49.4]
  reg [31:0] _RAND_23;
  reg [15:0] _T_83; // @[FIFO.scala 14:16:@50.4]
  reg [31:0] _RAND_24;
  reg [15:0] _T_86; // @[FIFO.scala 14:16:@51.4]
  reg [31:0] _RAND_25;
  reg [15:0] _T_89; // @[FIFO.scala 14:16:@52.4]
  reg [31:0] _RAND_26;
  reg [15:0] _T_92; // @[FIFO.scala 14:16:@53.4]
  reg [31:0] _RAND_27;
  reg [15:0] _T_95; // @[FIFO.scala 14:16:@54.4]
  reg [31:0] _RAND_28;
  reg [15:0] _T_98; // @[FIFO.scala 14:16:@55.4]
  reg [31:0] _RAND_29;
  reg [15:0] _T_101; // @[FIFO.scala 14:16:@56.4]
  reg [31:0] _RAND_30;
  reg [15:0] _T_104; // @[FIFO.scala 14:16:@57.4]
  reg [31:0] _RAND_31;
  reg [15:0] _T_107; // @[FIFO.scala 14:16:@58.4]
  reg [31:0] _RAND_32;
  reg [15:0] _T_110; // @[FIFO.scala 14:16:@59.4]
  reg [31:0] _RAND_33;
  reg [15:0] _T_113; // @[FIFO.scala 14:16:@60.4]
  reg [31:0] _RAND_34;
  reg [15:0] _T_116; // @[FIFO.scala 14:16:@61.4]
  reg [31:0] _RAND_35;
  reg [15:0] _T_119; // @[FIFO.scala 14:16:@62.4]
  reg [31:0] _RAND_36;
  reg [15:0] _T_122; // @[FIFO.scala 14:16:@63.4]
  reg [31:0] _RAND_37;
  reg [15:0] _T_125; // @[FIFO.scala 14:16:@64.4]
  reg [31:0] _RAND_38;
  reg [15:0] _T_128; // @[FIFO.scala 14:16:@65.4]
  reg [31:0] _RAND_39;
  reg [15:0] _T_131; // @[FIFO.scala 14:16:@66.4]
  reg [31:0] _RAND_40;
  reg [15:0] _T_134; // @[FIFO.scala 14:16:@67.4]
  reg [31:0] _RAND_41;
  reg [15:0] _T_137; // @[FIFO.scala 14:16:@68.4]
  reg [31:0] _RAND_42;
  reg [15:0] _T_140; // @[FIFO.scala 14:16:@69.4]
  reg [31:0] _RAND_43;
  reg [15:0] _T_143; // @[FIFO.scala 14:16:@70.4]
  reg [31:0] _RAND_44;
  reg [15:0] _T_146; // @[FIFO.scala 14:16:@71.4]
  reg [31:0] _RAND_45;
  reg [15:0] _T_149; // @[FIFO.scala 14:16:@72.4]
  reg [31:0] _RAND_46;
  reg [15:0] _T_152; // @[FIFO.scala 14:16:@73.4]
  reg [31:0] _RAND_47;
  reg [15:0] _T_155; // @[FIFO.scala 14:16:@74.4]
  reg [31:0] _RAND_48;
  reg [15:0] _T_158; // @[FIFO.scala 14:16:@75.4]
  reg [31:0] _RAND_49;
  reg [15:0] _T_161; // @[FIFO.scala 14:16:@76.4]
  reg [31:0] _RAND_50;
  reg [15:0] _T_164; // @[FIFO.scala 14:16:@77.4]
  reg [31:0] _RAND_51;
  reg [15:0] _T_167; // @[FIFO.scala 14:16:@78.4]
  reg [31:0] _RAND_52;
  reg [15:0] _T_170; // @[FIFO.scala 14:16:@79.4]
  reg [31:0] _RAND_53;
  reg [15:0] _T_173; // @[FIFO.scala 14:16:@80.4]
  reg [31:0] _RAND_54;
  reg [15:0] _T_176; // @[FIFO.scala 14:16:@81.4]
  reg [31:0] _RAND_55;
  reg [15:0] _T_179; // @[FIFO.scala 14:16:@82.4]
  reg [31:0] _RAND_56;
  reg [15:0] _T_182; // @[FIFO.scala 14:16:@83.4]
  reg [31:0] _RAND_57;
  reg [15:0] _T_185; // @[FIFO.scala 14:16:@84.4]
  reg [31:0] _RAND_58;
  reg [15:0] _T_188; // @[FIFO.scala 14:16:@85.4]
  reg [31:0] _RAND_59;
  reg [15:0] _T_191; // @[FIFO.scala 14:16:@86.4]
  reg [31:0] _RAND_60;
  reg [15:0] _T_194; // @[FIFO.scala 14:16:@87.4]
  reg [31:0] _RAND_61;
  reg [15:0] _T_197; // @[FIFO.scala 14:16:@88.4]
  reg [31:0] _RAND_62;
  reg [15:0] _T_200; // @[FIFO.scala 14:16:@89.4]
  reg [31:0] _RAND_63;
  reg [15:0] _T_203; // @[FIFO.scala 14:16:@90.4]
  reg [31:0] _RAND_64;
  reg [15:0] _T_206; // @[FIFO.scala 14:16:@91.4]
  reg [31:0] _RAND_65;
  reg [15:0] _T_209; // @[FIFO.scala 14:16:@92.4]
  reg [31:0] _RAND_66;
  reg [15:0] _T_212; // @[FIFO.scala 14:16:@93.4]
  reg [31:0] _RAND_67;
  reg [15:0] _T_215; // @[FIFO.scala 14:16:@94.4]
  reg [31:0] _RAND_68;
  reg [15:0] _T_218; // @[FIFO.scala 14:16:@95.4]
  reg [31:0] _RAND_69;
  reg [15:0] _T_221; // @[FIFO.scala 14:16:@96.4]
  reg [31:0] _RAND_70;
  reg [15:0] _T_224; // @[FIFO.scala 14:16:@97.4]
  reg [31:0] _RAND_71;
  reg [15:0] _T_227; // @[FIFO.scala 14:16:@98.4]
  reg [31:0] _RAND_72;
  reg [15:0] _T_230; // @[FIFO.scala 14:16:@99.4]
  reg [31:0] _RAND_73;
  reg [15:0] _T_233; // @[FIFO.scala 14:16:@100.4]
  reg [31:0] _RAND_74;
  reg [15:0] _T_236; // @[FIFO.scala 14:16:@101.4]
  reg [31:0] _RAND_75;
  reg [15:0] _T_239; // @[FIFO.scala 14:16:@102.4]
  reg [31:0] _RAND_76;
  reg [15:0] _T_242; // @[FIFO.scala 14:16:@103.4]
  reg [31:0] _RAND_77;
  reg [15:0] _T_245; // @[FIFO.scala 14:16:@104.4]
  reg [31:0] _RAND_78;
  reg [15:0] _T_248; // @[FIFO.scala 14:16:@105.4]
  reg [31:0] _RAND_79;
  reg [15:0] _T_251; // @[FIFO.scala 14:16:@106.4]
  reg [31:0] _RAND_80;
  reg [15:0] _T_254; // @[FIFO.scala 14:16:@107.4]
  reg [31:0] _RAND_81;
  reg [15:0] _T_257; // @[FIFO.scala 14:16:@108.4]
  reg [31:0] _RAND_82;
  reg [15:0] _T_260; // @[FIFO.scala 14:16:@109.4]
  reg [31:0] _RAND_83;
  reg [15:0] _T_263; // @[FIFO.scala 14:16:@110.4]
  reg [31:0] _RAND_84;
  reg [15:0] _T_266; // @[FIFO.scala 14:16:@111.4]
  reg [31:0] _RAND_85;
  reg [15:0] _T_269; // @[FIFO.scala 14:16:@112.4]
  reg [31:0] _RAND_86;
  reg [15:0] _T_272; // @[FIFO.scala 14:16:@113.4]
  reg [31:0] _RAND_87;
  reg [15:0] _T_275; // @[FIFO.scala 14:16:@114.4]
  reg [31:0] _RAND_88;
  reg [15:0] _T_278; // @[FIFO.scala 14:16:@115.4]
  reg [31:0] _RAND_89;
  reg [15:0] _T_281; // @[FIFO.scala 14:16:@116.4]
  reg [31:0] _RAND_90;
  reg [15:0] _T_284; // @[FIFO.scala 14:16:@117.4]
  reg [31:0] _RAND_91;
  reg [15:0] _T_287; // @[FIFO.scala 14:16:@118.4]
  reg [31:0] _RAND_92;
  reg [15:0] _T_290; // @[FIFO.scala 14:16:@119.4]
  reg [31:0] _RAND_93;
  reg [15:0] _T_293; // @[FIFO.scala 14:16:@120.4]
  reg [31:0] _RAND_94;
  reg [15:0] _T_296; // @[FIFO.scala 14:16:@121.4]
  reg [31:0] _RAND_95;
  reg [15:0] _T_299; // @[FIFO.scala 14:16:@122.4]
  reg [31:0] _RAND_96;
  reg [15:0] _T_302; // @[FIFO.scala 14:16:@123.4]
  reg [31:0] _RAND_97;
  reg [15:0] _T_305; // @[FIFO.scala 14:16:@124.4]
  reg [31:0] _RAND_98;
  reg [15:0] _T_308; // @[FIFO.scala 14:16:@125.4]
  reg [31:0] _RAND_99;
  reg [15:0] _T_311; // @[FIFO.scala 14:16:@126.4]
  reg [31:0] _RAND_100;
  reg [15:0] _T_314; // @[FIFO.scala 14:16:@127.4]
  reg [31:0] _RAND_101;
  reg [15:0] _T_317; // @[FIFO.scala 14:16:@128.4]
  reg [31:0] _RAND_102;
  reg [15:0] _T_320; // @[FIFO.scala 14:16:@129.4]
  reg [31:0] _RAND_103;
  reg [15:0] _T_323; // @[FIFO.scala 14:16:@130.4]
  reg [31:0] _RAND_104;
  reg [15:0] _T_326; // @[FIFO.scala 14:16:@131.4]
  reg [31:0] _RAND_105;
  reg [15:0] _T_329; // @[FIFO.scala 14:16:@132.4]
  reg [31:0] _RAND_106;
  reg [15:0] _T_332; // @[FIFO.scala 14:16:@133.4]
  reg [31:0] _RAND_107;
  reg [15:0] _T_335; // @[FIFO.scala 14:16:@134.4]
  reg [31:0] _RAND_108;
  reg [15:0] _T_338; // @[FIFO.scala 14:16:@135.4]
  reg [31:0] _RAND_109;
  reg [15:0] _T_341; // @[FIFO.scala 14:16:@136.4]
  reg [31:0] _RAND_110;
  reg [15:0] _T_344; // @[FIFO.scala 14:16:@137.4]
  reg [31:0] _RAND_111;
  reg [15:0] _T_347; // @[FIFO.scala 14:16:@138.4]
  reg [31:0] _RAND_112;
  reg [15:0] _T_350; // @[FIFO.scala 14:16:@139.4]
  reg [31:0] _RAND_113;
  reg [15:0] _T_353; // @[FIFO.scala 14:16:@140.4]
  reg [31:0] _RAND_114;
  reg [15:0] _T_356; // @[FIFO.scala 14:16:@141.4]
  reg [31:0] _RAND_115;
  reg [15:0] _T_359; // @[FIFO.scala 14:16:@142.4]
  reg [31:0] _RAND_116;
  reg [15:0] _T_362; // @[FIFO.scala 14:16:@143.4]
  reg [31:0] _RAND_117;
  reg [15:0] _T_365; // @[FIFO.scala 14:16:@144.4]
  reg [31:0] _RAND_118;
  reg [15:0] _T_368; // @[FIFO.scala 14:16:@145.4]
  reg [31:0] _RAND_119;
  reg [15:0] _T_371; // @[FIFO.scala 14:16:@146.4]
  reg [31:0] _RAND_120;
  reg [15:0] _T_374; // @[FIFO.scala 14:16:@147.4]
  reg [31:0] _RAND_121;
  reg [15:0] _T_377; // @[FIFO.scala 14:16:@148.4]
  reg [31:0] _RAND_122;
  reg [15:0] _T_380; // @[FIFO.scala 14:16:@149.4]
  reg [31:0] _RAND_123;
  reg [15:0] _T_383; // @[FIFO.scala 14:16:@150.4]
  reg [31:0] _RAND_124;
  reg [15:0] _T_386; // @[FIFO.scala 14:16:@151.4]
  reg [31:0] _RAND_125;
  reg [15:0] _T_389; // @[FIFO.scala 14:16:@152.4]
  reg [31:0] _RAND_126;
  reg [15:0] _T_392; // @[FIFO.scala 14:16:@153.4]
  reg [31:0] _RAND_127;
  reg [15:0] _T_395; // @[FIFO.scala 14:16:@154.4]
  reg [31:0] _RAND_128;
  reg [15:0] _T_398; // @[FIFO.scala 14:16:@155.4]
  reg [31:0] _RAND_129;
  reg [15:0] _T_401; // @[FIFO.scala 14:16:@156.4]
  reg [31:0] _RAND_130;
  reg [15:0] _T_404; // @[FIFO.scala 14:16:@157.4]
  reg [31:0] _RAND_131;
  reg [15:0] _T_407; // @[FIFO.scala 14:16:@158.4]
  reg [31:0] _RAND_132;
  reg [15:0] _T_410; // @[FIFO.scala 14:16:@159.4]
  reg [31:0] _RAND_133;
  reg [15:0] _T_413; // @[FIFO.scala 14:16:@160.4]
  reg [31:0] _RAND_134;
  reg [15:0] _T_416; // @[FIFO.scala 14:16:@161.4]
  reg [31:0] _RAND_135;
  reg [15:0] _T_419; // @[FIFO.scala 14:16:@162.4]
  reg [31:0] _RAND_136;
  reg [15:0] _T_422; // @[FIFO.scala 14:16:@163.4]
  reg [31:0] _RAND_137;
  reg [15:0] _T_425; // @[FIFO.scala 14:16:@164.4]
  reg [31:0] _RAND_138;
  reg [15:0] _T_428; // @[FIFO.scala 14:16:@165.4]
  reg [31:0] _RAND_139;
  reg [15:0] _T_431; // @[FIFO.scala 14:16:@166.4]
  reg [31:0] _RAND_140;
  reg [15:0] _T_434; // @[FIFO.scala 14:16:@167.4]
  reg [31:0] _RAND_141;
  reg [15:0] _T_437; // @[FIFO.scala 14:16:@168.4]
  reg [31:0] _RAND_142;
  reg [15:0] _T_440; // @[FIFO.scala 14:16:@169.4]
  reg [31:0] _RAND_143;
  reg [15:0] _T_443; // @[FIFO.scala 14:16:@170.4]
  reg [31:0] _RAND_144;
  reg [15:0] _T_446; // @[FIFO.scala 14:16:@171.4]
  reg [31:0] _RAND_145;
  reg [15:0] _T_449; // @[FIFO.scala 14:16:@172.4]
  reg [31:0] _RAND_146;
  reg [15:0] _T_452; // @[FIFO.scala 14:16:@173.4]
  reg [31:0] _RAND_147;
  reg [15:0] _T_455; // @[FIFO.scala 14:16:@174.4]
  reg [31:0] _RAND_148;
  reg [15:0] _T_458; // @[FIFO.scala 14:16:@175.4]
  reg [31:0] _RAND_149;
  reg [15:0] _T_461; // @[FIFO.scala 14:16:@176.4]
  reg [31:0] _RAND_150;
  reg [15:0] _T_464; // @[FIFO.scala 14:16:@177.4]
  reg [31:0] _RAND_151;
  reg [15:0] _T_467; // @[FIFO.scala 14:16:@178.4]
  reg [31:0] _RAND_152;
  reg [15:0] _T_470; // @[FIFO.scala 14:16:@179.4]
  reg [31:0] _RAND_153;
  reg [15:0] _T_473; // @[FIFO.scala 14:16:@180.4]
  reg [31:0] _RAND_154;
  reg [15:0] _T_476; // @[FIFO.scala 14:16:@181.4]
  reg [31:0] _RAND_155;
  reg [15:0] _T_479; // @[FIFO.scala 14:16:@182.4]
  reg [31:0] _RAND_156;
  reg [15:0] _T_482; // @[FIFO.scala 14:16:@183.4]
  reg [31:0] _RAND_157;
  reg [15:0] _T_485; // @[FIFO.scala 14:16:@184.4]
  reg [31:0] _RAND_158;
  reg [15:0] _T_488; // @[FIFO.scala 14:16:@185.4]
  reg [31:0] _RAND_159;
  reg [15:0] _T_491; // @[FIFO.scala 14:16:@186.4]
  reg [31:0] _RAND_160;
  reg [15:0] _T_494; // @[FIFO.scala 14:16:@187.4]
  reg [31:0] _RAND_161;
  reg [15:0] _T_497; // @[FIFO.scala 14:16:@188.4]
  reg [31:0] _RAND_162;
  reg [15:0] _T_500; // @[FIFO.scala 14:16:@189.4]
  reg [31:0] _RAND_163;
  reg [15:0] _T_503; // @[FIFO.scala 14:16:@190.4]
  reg [31:0] _RAND_164;
  reg [15:0] _T_506; // @[FIFO.scala 14:16:@191.4]
  reg [31:0] _RAND_165;
  reg [15:0] _T_509; // @[FIFO.scala 14:16:@192.4]
  reg [31:0] _RAND_166;
  reg [15:0] _T_512; // @[FIFO.scala 14:16:@193.4]
  reg [31:0] _RAND_167;
  reg [15:0] _T_515; // @[FIFO.scala 14:16:@194.4]
  reg [31:0] _RAND_168;
  reg [15:0] _T_518; // @[FIFO.scala 14:16:@195.4]
  reg [31:0] _RAND_169;
  reg [15:0] _T_521; // @[FIFO.scala 14:16:@196.4]
  reg [31:0] _RAND_170;
  reg [15:0] _T_524; // @[FIFO.scala 14:16:@197.4]
  reg [31:0] _RAND_171;
  reg [15:0] _T_527; // @[FIFO.scala 14:16:@198.4]
  reg [31:0] _RAND_172;
  reg [15:0] _T_530; // @[FIFO.scala 14:16:@199.4]
  reg [31:0] _RAND_173;
  reg [15:0] _T_533; // @[FIFO.scala 14:16:@200.4]
  reg [31:0] _RAND_174;
  reg [15:0] _T_536; // @[FIFO.scala 14:16:@201.4]
  reg [31:0] _RAND_175;
  reg [15:0] _T_539; // @[FIFO.scala 14:16:@202.4]
  reg [31:0] _RAND_176;
  reg [15:0] _T_542; // @[FIFO.scala 14:16:@203.4]
  reg [31:0] _RAND_177;
  reg [15:0] _T_545; // @[FIFO.scala 14:16:@204.4]
  reg [31:0] _RAND_178;
  reg [15:0] _T_548; // @[FIFO.scala 14:16:@205.4]
  reg [31:0] _RAND_179;
  reg [15:0] _T_551; // @[FIFO.scala 14:16:@206.4]
  reg [31:0] _RAND_180;
  reg [15:0] _T_554; // @[FIFO.scala 14:16:@207.4]
  reg [31:0] _RAND_181;
  reg [15:0] _T_557; // @[FIFO.scala 14:16:@208.4]
  reg [31:0] _RAND_182;
  reg [15:0] _T_560; // @[FIFO.scala 14:16:@209.4]
  reg [31:0] _RAND_183;
  reg [15:0] _T_563; // @[FIFO.scala 14:16:@210.4]
  reg [31:0] _RAND_184;
  reg [15:0] _T_566; // @[FIFO.scala 14:16:@211.4]
  reg [31:0] _RAND_185;
  reg [15:0] _T_569; // @[FIFO.scala 14:16:@212.4]
  reg [31:0] _RAND_186;
  reg [15:0] _T_572; // @[FIFO.scala 14:16:@213.4]
  reg [31:0] _RAND_187;
  reg [15:0] _T_575; // @[FIFO.scala 14:16:@214.4]
  reg [31:0] _RAND_188;
  reg [15:0] _T_578; // @[FIFO.scala 14:16:@215.4]
  reg [31:0] _RAND_189;
  reg [15:0] _T_581; // @[FIFO.scala 14:16:@216.4]
  reg [31:0] _RAND_190;
  reg [15:0] _T_584; // @[FIFO.scala 14:16:@217.4]
  reg [31:0] _RAND_191;
  reg [15:0] _T_587; // @[FIFO.scala 14:16:@218.4]
  reg [31:0] _RAND_192;
  reg [15:0] _T_590; // @[FIFO.scala 14:16:@219.4]
  reg [31:0] _RAND_193;
  reg [15:0] _T_593; // @[FIFO.scala 14:16:@220.4]
  reg [31:0] _RAND_194;
  reg [15:0] _T_596; // @[FIFO.scala 14:16:@221.4]
  reg [31:0] _RAND_195;
  reg [15:0] _T_599; // @[FIFO.scala 14:16:@222.4]
  reg [31:0] _RAND_196;
  reg [15:0] _T_602; // @[FIFO.scala 14:16:@223.4]
  reg [31:0] _RAND_197;
  reg [15:0] _T_605; // @[FIFO.scala 14:16:@224.4]
  reg [31:0] _RAND_198;
  reg [15:0] _T_608; // @[FIFO.scala 14:16:@225.4]
  reg [31:0] _RAND_199;
  reg [15:0] _T_611; // @[FIFO.scala 14:16:@226.4]
  reg [31:0] _RAND_200;
  reg [15:0] _T_614; // @[FIFO.scala 14:16:@227.4]
  reg [31:0] _RAND_201;
  reg [15:0] _T_617; // @[FIFO.scala 14:16:@228.4]
  reg [31:0] _RAND_202;
  reg [15:0] _T_620; // @[FIFO.scala 14:16:@229.4]
  reg [31:0] _RAND_203;
  reg [15:0] _T_623; // @[FIFO.scala 14:16:@230.4]
  reg [31:0] _RAND_204;
  reg [15:0] _T_626; // @[FIFO.scala 14:16:@231.4]
  reg [31:0] _RAND_205;
  reg [15:0] _T_629; // @[FIFO.scala 14:16:@232.4]
  reg [31:0] _RAND_206;
  reg [15:0] _T_632; // @[FIFO.scala 14:16:@233.4]
  reg [31:0] _RAND_207;
  reg [15:0] _T_635; // @[FIFO.scala 14:16:@234.4]
  reg [31:0] _RAND_208;
  reg [15:0] _T_638; // @[FIFO.scala 14:16:@235.4]
  reg [31:0] _RAND_209;
  reg [15:0] _T_641; // @[FIFO.scala 14:16:@236.4]
  reg [31:0] _RAND_210;
  reg [15:0] _T_644; // @[FIFO.scala 14:16:@237.4]
  reg [31:0] _RAND_211;
  reg [15:0] _T_647; // @[FIFO.scala 14:16:@238.4]
  reg [31:0] _RAND_212;
  reg [15:0] _T_650; // @[FIFO.scala 14:16:@239.4]
  reg [31:0] _RAND_213;
  reg [15:0] _T_653; // @[FIFO.scala 14:16:@240.4]
  reg [31:0] _RAND_214;
  reg [15:0] _T_656; // @[FIFO.scala 14:16:@241.4]
  reg [31:0] _RAND_215;
  reg [15:0] _T_659; // @[FIFO.scala 14:16:@242.4]
  reg [31:0] _RAND_216;
  reg [15:0] _T_662; // @[FIFO.scala 14:16:@243.4]
  reg [31:0] _RAND_217;
  reg [15:0] _T_665; // @[FIFO.scala 14:16:@244.4]
  reg [31:0] _RAND_218;
  reg [15:0] _T_668; // @[FIFO.scala 14:16:@245.4]
  reg [31:0] _RAND_219;
  reg [15:0] _T_671; // @[FIFO.scala 14:16:@246.4]
  reg [31:0] _RAND_220;
  reg [15:0] _T_674; // @[FIFO.scala 14:16:@247.4]
  reg [31:0] _RAND_221;
  reg [15:0] _T_677; // @[FIFO.scala 14:16:@248.4]
  reg [31:0] _RAND_222;
  reg [15:0] _T_680; // @[FIFO.scala 14:16:@249.4]
  reg [31:0] _RAND_223;
  reg [15:0] _T_683; // @[FIFO.scala 14:16:@250.4]
  reg [31:0] _RAND_224;
  reg [15:0] _T_686; // @[FIFO.scala 14:16:@251.4]
  reg [31:0] _RAND_225;
  reg [15:0] _T_689; // @[FIFO.scala 14:16:@252.4]
  reg [31:0] _RAND_226;
  reg [15:0] _T_692; // @[FIFO.scala 14:16:@253.4]
  reg [31:0] _RAND_227;
  reg [15:0] _T_695; // @[FIFO.scala 14:16:@254.4]
  reg [31:0] _RAND_228;
  reg [15:0] _T_698; // @[FIFO.scala 14:16:@255.4]
  reg [31:0] _RAND_229;
  reg [15:0] _T_701; // @[FIFO.scala 14:16:@256.4]
  reg [31:0] _RAND_230;
  reg [15:0] _T_704; // @[FIFO.scala 14:16:@257.4]
  reg [31:0] _RAND_231;
  reg [15:0] _T_707; // @[FIFO.scala 14:16:@258.4]
  reg [31:0] _RAND_232;
  reg [15:0] _T_710; // @[FIFO.scala 14:16:@259.4]
  reg [31:0] _RAND_233;
  reg [15:0] _T_713; // @[FIFO.scala 14:16:@260.4]
  reg [31:0] _RAND_234;
  reg [15:0] _T_716; // @[FIFO.scala 14:16:@261.4]
  reg [31:0] _RAND_235;
  reg [15:0] _T_719; // @[FIFO.scala 14:16:@262.4]
  reg [31:0] _RAND_236;
  reg [15:0] _T_722; // @[FIFO.scala 14:16:@263.4]
  reg [31:0] _RAND_237;
  reg [15:0] _T_725; // @[FIFO.scala 14:16:@264.4]
  reg [31:0] _RAND_238;
  reg [15:0] _T_728; // @[FIFO.scala 14:16:@265.4]
  reg [31:0] _RAND_239;
  reg [15:0] _T_731; // @[FIFO.scala 14:16:@266.4]
  reg [31:0] _RAND_240;
  reg [15:0] _T_734; // @[FIFO.scala 14:16:@267.4]
  reg [31:0] _RAND_241;
  reg [15:0] _T_737; // @[FIFO.scala 14:16:@268.4]
  reg [31:0] _RAND_242;
  reg [15:0] _T_740; // @[FIFO.scala 14:16:@269.4]
  reg [31:0] _RAND_243;
  reg [15:0] _T_743; // @[FIFO.scala 14:16:@270.4]
  reg [31:0] _RAND_244;
  reg [15:0] _T_746; // @[FIFO.scala 14:16:@271.4]
  reg [31:0] _RAND_245;
  reg [15:0] _T_749; // @[FIFO.scala 14:16:@272.4]
  reg [31:0] _RAND_246;
  reg [15:0] _T_752; // @[FIFO.scala 14:16:@273.4]
  reg [31:0] _RAND_247;
  reg [15:0] _T_755; // @[FIFO.scala 14:16:@274.4]
  reg [31:0] _RAND_248;
  reg [15:0] _T_758; // @[FIFO.scala 14:16:@275.4]
  reg [31:0] _RAND_249;
  reg [15:0] _T_761; // @[FIFO.scala 14:16:@276.4]
  reg [31:0] _RAND_250;
  reg [15:0] _T_764; // @[FIFO.scala 14:16:@277.4]
  reg [31:0] _RAND_251;
  reg [15:0] _T_767; // @[FIFO.scala 14:16:@278.4]
  reg [31:0] _RAND_252;
  reg [15:0] _T_770; // @[FIFO.scala 14:16:@279.4]
  reg [31:0] _RAND_253;
  reg [15:0] _T_773; // @[FIFO.scala 14:16:@280.4]
  reg [31:0] _RAND_254;
  reg [15:0] _T_776; // @[FIFO.scala 14:16:@281.4]
  reg [31:0] _RAND_255;
  reg [15:0] _T_779; // @[FIFO.scala 14:16:@282.4]
  reg [31:0] _RAND_256;
  reg [15:0] _T_782; // @[FIFO.scala 14:16:@283.4]
  reg [31:0] _RAND_257;
  reg [15:0] _T_785; // @[FIFO.scala 14:16:@284.4]
  reg [31:0] _RAND_258;
  reg [15:0] _T_788; // @[FIFO.scala 14:16:@285.4]
  reg [31:0] _RAND_259;
  reg [15:0] _T_791; // @[FIFO.scala 14:16:@286.4]
  reg [31:0] _RAND_260;
  reg [15:0] _T_794; // @[FIFO.scala 14:16:@287.4]
  reg [31:0] _RAND_261;
  reg [15:0] _T_797; // @[FIFO.scala 14:16:@288.4]
  reg [31:0] _RAND_262;
  reg [15:0] _T_800; // @[FIFO.scala 14:16:@289.4]
  reg [31:0] _RAND_263;
  reg [15:0] _T_803; // @[FIFO.scala 14:16:@290.4]
  reg [31:0] _RAND_264;
  reg [15:0] _T_806; // @[FIFO.scala 14:16:@291.4]
  reg [31:0] _RAND_265;
  reg [15:0] _T_809; // @[FIFO.scala 14:16:@292.4]
  reg [31:0] _RAND_266;
  reg [15:0] _T_812; // @[FIFO.scala 14:16:@293.4]
  reg [31:0] _RAND_267;
  reg [15:0] _T_815; // @[FIFO.scala 14:16:@294.4]
  reg [31:0] _RAND_268;
  reg [15:0] _T_818; // @[FIFO.scala 14:16:@295.4]
  reg [31:0] _RAND_269;
  reg [15:0] _T_821; // @[FIFO.scala 14:16:@296.4]
  reg [31:0] _RAND_270;
  reg [15:0] _T_824; // @[FIFO.scala 14:16:@297.4]
  reg [31:0] _RAND_271;
  reg [15:0] _T_827; // @[FIFO.scala 14:16:@298.4]
  reg [31:0] _RAND_272;
  reg [15:0] _T_830; // @[FIFO.scala 14:16:@299.4]
  reg [31:0] _RAND_273;
  reg [15:0] _T_833; // @[FIFO.scala 14:16:@300.4]
  reg [31:0] _RAND_274;
  reg [15:0] _T_836; // @[FIFO.scala 14:16:@301.4]
  reg [31:0] _RAND_275;
  reg [15:0] _T_839; // @[FIFO.scala 14:16:@302.4]
  reg [31:0] _RAND_276;
  reg [15:0] _T_842; // @[FIFO.scala 14:16:@303.4]
  reg [31:0] _RAND_277;
  reg [15:0] _T_845; // @[FIFO.scala 14:16:@304.4]
  reg [31:0] _RAND_278;
  reg [15:0] _T_848; // @[FIFO.scala 14:16:@305.4]
  reg [31:0] _RAND_279;
  reg [15:0] _T_851; // @[FIFO.scala 14:16:@306.4]
  reg [31:0] _RAND_280;
  reg [15:0] _T_854; // @[FIFO.scala 14:16:@307.4]
  reg [31:0] _RAND_281;
  reg [15:0] _T_857; // @[FIFO.scala 14:16:@308.4]
  reg [31:0] _RAND_282;
  reg [15:0] _T_860; // @[FIFO.scala 14:16:@309.4]
  reg [31:0] _RAND_283;
  reg [15:0] _T_863; // @[FIFO.scala 14:16:@310.4]
  reg [31:0] _RAND_284;
  reg [15:0] _T_866; // @[FIFO.scala 14:16:@311.4]
  reg [31:0] _RAND_285;
  reg [15:0] _T_869; // @[FIFO.scala 14:16:@312.4]
  reg [31:0] _RAND_286;
  reg [15:0] _T_872; // @[FIFO.scala 14:16:@313.4]
  reg [31:0] _RAND_287;
  reg [15:0] _T_875; // @[FIFO.scala 14:16:@314.4]
  reg [31:0] _RAND_288;
  reg [15:0] _T_878; // @[FIFO.scala 14:16:@315.4]
  reg [31:0] _RAND_289;
  reg [15:0] _T_881; // @[FIFO.scala 14:16:@316.4]
  reg [31:0] _RAND_290;
  reg [15:0] _T_884; // @[FIFO.scala 14:16:@317.4]
  reg [31:0] _RAND_291;
  reg [15:0] _T_887; // @[FIFO.scala 14:16:@318.4]
  reg [31:0] _RAND_292;
  reg [15:0] _T_890; // @[FIFO.scala 14:16:@319.4]
  reg [31:0] _RAND_293;
  reg [15:0] _T_893; // @[FIFO.scala 14:16:@320.4]
  reg [31:0] _RAND_294;
  reg [15:0] _T_896; // @[FIFO.scala 14:16:@321.4]
  reg [31:0] _RAND_295;
  reg [15:0] _T_899; // @[FIFO.scala 14:16:@322.4]
  reg [31:0] _RAND_296;
  reg [15:0] _T_902; // @[FIFO.scala 14:16:@323.4]
  reg [31:0] _RAND_297;
  reg [15:0] _T_905; // @[FIFO.scala 14:16:@324.4]
  reg [31:0] _RAND_298;
  reg [15:0] _T_908; // @[FIFO.scala 14:16:@325.4]
  reg [31:0] _RAND_299;
  reg [15:0] _T_911; // @[FIFO.scala 14:16:@326.4]
  reg [31:0] _RAND_300;
  reg [15:0] _T_914; // @[FIFO.scala 14:16:@327.4]
  reg [31:0] _RAND_301;
  reg [15:0] _T_917; // @[FIFO.scala 14:16:@328.4]
  reg [31:0] _RAND_302;
  reg [15:0] _T_920; // @[FIFO.scala 14:16:@329.4]
  reg [31:0] _RAND_303;
  reg [15:0] _T_923; // @[FIFO.scala 14:16:@330.4]
  reg [31:0] _RAND_304;
  reg [15:0] _T_926; // @[FIFO.scala 14:16:@331.4]
  reg [31:0] _RAND_305;
  reg [15:0] _T_929; // @[FIFO.scala 14:16:@332.4]
  reg [31:0] _RAND_306;
  reg [15:0] _T_932; // @[FIFO.scala 14:16:@333.4]
  reg [31:0] _RAND_307;
  reg [15:0] _T_935; // @[FIFO.scala 14:16:@334.4]
  reg [31:0] _RAND_308;
  reg [15:0] _T_938; // @[FIFO.scala 14:16:@335.4]
  reg [31:0] _RAND_309;
  reg [15:0] _T_941; // @[FIFO.scala 14:16:@336.4]
  reg [31:0] _RAND_310;
  reg [15:0] _T_944; // @[FIFO.scala 14:16:@337.4]
  reg [31:0] _RAND_311;
  reg [15:0] _T_947; // @[FIFO.scala 14:16:@338.4]
  reg [31:0] _RAND_312;
  reg [15:0] _T_950; // @[FIFO.scala 14:16:@339.4]
  reg [31:0] _RAND_313;
  reg [15:0] _T_953; // @[FIFO.scala 14:16:@340.4]
  reg [31:0] _RAND_314;
  reg [15:0] _T_956; // @[FIFO.scala 14:16:@341.4]
  reg [31:0] _RAND_315;
  reg [15:0] _T_959; // @[FIFO.scala 14:16:@342.4]
  reg [31:0] _RAND_316;
  assign io_dataOut = _T_959; // @[FIFO.scala 22:14:@659.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_11 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_14 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_17 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_20 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_23 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_26 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_29 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_32 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_35 = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_38 = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_41 = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_44 = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_47 = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_50 = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_53 = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_56 = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_59 = _RAND_16[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_62 = _RAND_17[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_65 = _RAND_18[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_68 = _RAND_19[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_71 = _RAND_20[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_74 = _RAND_21[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_77 = _RAND_22[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_80 = _RAND_23[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_83 = _RAND_24[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_86 = _RAND_25[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_89 = _RAND_26[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_92 = _RAND_27[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_95 = _RAND_28[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_98 = _RAND_29[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_101 = _RAND_30[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_104 = _RAND_31[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_107 = _RAND_32[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_110 = _RAND_33[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_113 = _RAND_34[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_116 = _RAND_35[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_119 = _RAND_36[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_122 = _RAND_37[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_125 = _RAND_38[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_128 = _RAND_39[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_131 = _RAND_40[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_134 = _RAND_41[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_137 = _RAND_42[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_140 = _RAND_43[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_143 = _RAND_44[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_146 = _RAND_45[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_149 = _RAND_46[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_152 = _RAND_47[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_155 = _RAND_48[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_158 = _RAND_49[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_161 = _RAND_50[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_164 = _RAND_51[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_167 = _RAND_52[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_170 = _RAND_53[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_173 = _RAND_54[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_176 = _RAND_55[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_179 = _RAND_56[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_182 = _RAND_57[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_185 = _RAND_58[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_188 = _RAND_59[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_191 = _RAND_60[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_194 = _RAND_61[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_197 = _RAND_62[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_200 = _RAND_63[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_203 = _RAND_64[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_206 = _RAND_65[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_209 = _RAND_66[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_212 = _RAND_67[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_215 = _RAND_68[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_218 = _RAND_69[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_221 = _RAND_70[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_224 = _RAND_71[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_227 = _RAND_72[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_230 = _RAND_73[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_233 = _RAND_74[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_236 = _RAND_75[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_239 = _RAND_76[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_242 = _RAND_77[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_245 = _RAND_78[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_248 = _RAND_79[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_251 = _RAND_80[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_254 = _RAND_81[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_257 = _RAND_82[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_260 = _RAND_83[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_263 = _RAND_84[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_266 = _RAND_85[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_269 = _RAND_86[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_272 = _RAND_87[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_275 = _RAND_88[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_278 = _RAND_89[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_281 = _RAND_90[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_284 = _RAND_91[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_287 = _RAND_92[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_290 = _RAND_93[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_293 = _RAND_94[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_296 = _RAND_95[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_299 = _RAND_96[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_302 = _RAND_97[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_305 = _RAND_98[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_308 = _RAND_99[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_311 = _RAND_100[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_314 = _RAND_101[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_317 = _RAND_102[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_320 = _RAND_103[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_323 = _RAND_104[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_326 = _RAND_105[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_329 = _RAND_106[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_332 = _RAND_107[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_335 = _RAND_108[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_338 = _RAND_109[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_341 = _RAND_110[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_344 = _RAND_111[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_347 = _RAND_112[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_350 = _RAND_113[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_353 = _RAND_114[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_356 = _RAND_115[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_359 = _RAND_116[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_362 = _RAND_117[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_365 = _RAND_118[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_368 = _RAND_119[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_371 = _RAND_120[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_374 = _RAND_121[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_377 = _RAND_122[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_380 = _RAND_123[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_383 = _RAND_124[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T_386 = _RAND_125[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_389 = _RAND_126[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_392 = _RAND_127[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_395 = _RAND_128[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T_398 = _RAND_129[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _T_401 = _RAND_130[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _T_404 = _RAND_131[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _T_407 = _RAND_132[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _T_410 = _RAND_133[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _T_413 = _RAND_134[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _T_416 = _RAND_135[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _T_419 = _RAND_136[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _T_422 = _RAND_137[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _T_425 = _RAND_138[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _T_428 = _RAND_139[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _T_431 = _RAND_140[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _T_434 = _RAND_141[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _T_437 = _RAND_142[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _T_440 = _RAND_143[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _T_443 = _RAND_144[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _T_446 = _RAND_145[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _T_449 = _RAND_146[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  _T_452 = _RAND_147[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  _T_455 = _RAND_148[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  _T_458 = _RAND_149[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _T_461 = _RAND_150[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _T_464 = _RAND_151[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  _T_467 = _RAND_152[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _T_470 = _RAND_153[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _T_473 = _RAND_154[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _T_476 = _RAND_155[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _T_479 = _RAND_156[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _T_482 = _RAND_157[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _T_485 = _RAND_158[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _T_488 = _RAND_159[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _T_491 = _RAND_160[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _T_494 = _RAND_161[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _T_497 = _RAND_162[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _T_500 = _RAND_163[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _T_503 = _RAND_164[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _T_506 = _RAND_165[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _T_509 = _RAND_166[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _T_512 = _RAND_167[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _T_515 = _RAND_168[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _T_518 = _RAND_169[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _T_521 = _RAND_170[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _T_524 = _RAND_171[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _T_527 = _RAND_172[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _T_530 = _RAND_173[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _T_533 = _RAND_174[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _T_536 = _RAND_175[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _T_539 = _RAND_176[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _T_542 = _RAND_177[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _T_545 = _RAND_178[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _T_548 = _RAND_179[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  _T_551 = _RAND_180[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _T_554 = _RAND_181[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _T_557 = _RAND_182[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _T_560 = _RAND_183[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _T_563 = _RAND_184[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _T_566 = _RAND_185[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _T_569 = _RAND_186[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _T_572 = _RAND_187[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _T_575 = _RAND_188[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _T_578 = _RAND_189[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _T_581 = _RAND_190[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  _T_584 = _RAND_191[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  _T_587 = _RAND_192[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  _T_590 = _RAND_193[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _T_593 = _RAND_194[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _T_596 = _RAND_195[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _T_599 = _RAND_196[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  _T_602 = _RAND_197[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  _T_605 = _RAND_198[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  _T_608 = _RAND_199[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _T_611 = _RAND_200[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  _T_614 = _RAND_201[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  _T_617 = _RAND_202[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  _T_620 = _RAND_203[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  _T_623 = _RAND_204[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  _T_626 = _RAND_205[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  _T_629 = _RAND_206[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  _T_632 = _RAND_207[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  _T_635 = _RAND_208[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  _T_638 = _RAND_209[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  _T_641 = _RAND_210[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  _T_644 = _RAND_211[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  _T_647 = _RAND_212[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  _T_650 = _RAND_213[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  _T_653 = _RAND_214[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  _T_656 = _RAND_215[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  _T_659 = _RAND_216[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  _T_662 = _RAND_217[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  _T_665 = _RAND_218[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  _T_668 = _RAND_219[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  _T_671 = _RAND_220[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  _T_674 = _RAND_221[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  _T_677 = _RAND_222[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  _T_680 = _RAND_223[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  _T_683 = _RAND_224[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  _T_686 = _RAND_225[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  _T_689 = _RAND_226[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  _T_692 = _RAND_227[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  _T_695 = _RAND_228[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  _T_698 = _RAND_229[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  _T_701 = _RAND_230[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  _T_704 = _RAND_231[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  _T_707 = _RAND_232[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  _T_710 = _RAND_233[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  _T_713 = _RAND_234[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  _T_716 = _RAND_235[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  _T_719 = _RAND_236[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  _T_722 = _RAND_237[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  _T_725 = _RAND_238[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  _T_728 = _RAND_239[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  _T_731 = _RAND_240[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  _T_734 = _RAND_241[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  _T_737 = _RAND_242[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  _T_740 = _RAND_243[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  _T_743 = _RAND_244[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  _T_746 = _RAND_245[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  _T_749 = _RAND_246[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  _T_752 = _RAND_247[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  _T_755 = _RAND_248[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  _T_758 = _RAND_249[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  _T_761 = _RAND_250[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  _T_764 = _RAND_251[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  _T_767 = _RAND_252[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  _T_770 = _RAND_253[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  _T_773 = _RAND_254[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  _T_776 = _RAND_255[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  _T_779 = _RAND_256[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  _T_782 = _RAND_257[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  _T_785 = _RAND_258[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  _T_788 = _RAND_259[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  _T_791 = _RAND_260[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  _T_794 = _RAND_261[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  _T_797 = _RAND_262[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  _T_800 = _RAND_263[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  _T_803 = _RAND_264[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  _T_806 = _RAND_265[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  _T_809 = _RAND_266[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  _T_812 = _RAND_267[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  _T_815 = _RAND_268[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  _T_818 = _RAND_269[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  _T_821 = _RAND_270[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  _T_824 = _RAND_271[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  _T_827 = _RAND_272[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  _T_830 = _RAND_273[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  _T_833 = _RAND_274[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  _T_836 = _RAND_275[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  _T_839 = _RAND_276[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  _T_842 = _RAND_277[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  _T_845 = _RAND_278[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  _T_848 = _RAND_279[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  _T_851 = _RAND_280[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  _T_854 = _RAND_281[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  _T_857 = _RAND_282[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  _T_860 = _RAND_283[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  _T_863 = _RAND_284[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  _T_866 = _RAND_285[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  _T_869 = _RAND_286[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  _T_872 = _RAND_287[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  _T_875 = _RAND_288[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  _T_878 = _RAND_289[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  _T_881 = _RAND_290[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  _T_884 = _RAND_291[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  _T_887 = _RAND_292[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  _T_890 = _RAND_293[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  _T_893 = _RAND_294[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  _T_896 = _RAND_295[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  _T_899 = _RAND_296[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  _T_902 = _RAND_297[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  _T_905 = _RAND_298[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  _T_908 = _RAND_299[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  _T_911 = _RAND_300[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  _T_914 = _RAND_301[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  _T_917 = _RAND_302[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  _T_920 = _RAND_303[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  _T_923 = _RAND_304[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  _T_926 = _RAND_305[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  _T_929 = _RAND_306[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  _T_932 = _RAND_307[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  _T_935 = _RAND_308[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  _T_938 = _RAND_309[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  _T_941 = _RAND_310[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  _T_944 = _RAND_311[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  _T_947 = _RAND_312[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  _T_950 = _RAND_313[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  _T_953 = _RAND_314[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  _T_956 = _RAND_315[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  _T_959 = _RAND_316[15:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_11 <= 16'sh0;
    end else begin
      _T_11 <= io_dataIn;
    end
    if (reset) begin
      _T_14 <= 16'sh0;
    end else begin
      _T_14 <= _T_11;
    end
    if (reset) begin
      _T_17 <= 16'sh0;
    end else begin
      _T_17 <= _T_14;
    end
    if (reset) begin
      _T_20 <= 16'sh0;
    end else begin
      _T_20 <= _T_17;
    end
    if (reset) begin
      _T_23 <= 16'sh0;
    end else begin
      _T_23 <= _T_20;
    end
    if (reset) begin
      _T_26 <= 16'sh0;
    end else begin
      _T_26 <= _T_23;
    end
    if (reset) begin
      _T_29 <= 16'sh0;
    end else begin
      _T_29 <= _T_26;
    end
    if (reset) begin
      _T_32 <= 16'sh0;
    end else begin
      _T_32 <= _T_29;
    end
    if (reset) begin
      _T_35 <= 16'sh0;
    end else begin
      _T_35 <= _T_32;
    end
    if (reset) begin
      _T_38 <= 16'sh0;
    end else begin
      _T_38 <= _T_35;
    end
    if (reset) begin
      _T_41 <= 16'sh0;
    end else begin
      _T_41 <= _T_38;
    end
    if (reset) begin
      _T_44 <= 16'sh0;
    end else begin
      _T_44 <= _T_41;
    end
    if (reset) begin
      _T_47 <= 16'sh0;
    end else begin
      _T_47 <= _T_44;
    end
    if (reset) begin
      _T_50 <= 16'sh0;
    end else begin
      _T_50 <= _T_47;
    end
    if (reset) begin
      _T_53 <= 16'sh0;
    end else begin
      _T_53 <= _T_50;
    end
    if (reset) begin
      _T_56 <= 16'sh0;
    end else begin
      _T_56 <= _T_53;
    end
    if (reset) begin
      _T_59 <= 16'sh0;
    end else begin
      _T_59 <= _T_56;
    end
    if (reset) begin
      _T_62 <= 16'sh0;
    end else begin
      _T_62 <= _T_59;
    end
    if (reset) begin
      _T_65 <= 16'sh0;
    end else begin
      _T_65 <= _T_62;
    end
    if (reset) begin
      _T_68 <= 16'sh0;
    end else begin
      _T_68 <= _T_65;
    end
    if (reset) begin
      _T_71 <= 16'sh0;
    end else begin
      _T_71 <= _T_68;
    end
    if (reset) begin
      _T_74 <= 16'sh0;
    end else begin
      _T_74 <= _T_71;
    end
    if (reset) begin
      _T_77 <= 16'sh0;
    end else begin
      _T_77 <= _T_74;
    end
    if (reset) begin
      _T_80 <= 16'sh0;
    end else begin
      _T_80 <= _T_77;
    end
    if (reset) begin
      _T_83 <= 16'sh0;
    end else begin
      _T_83 <= _T_80;
    end
    if (reset) begin
      _T_86 <= 16'sh0;
    end else begin
      _T_86 <= _T_83;
    end
    if (reset) begin
      _T_89 <= 16'sh0;
    end else begin
      _T_89 <= _T_86;
    end
    if (reset) begin
      _T_92 <= 16'sh0;
    end else begin
      _T_92 <= _T_89;
    end
    if (reset) begin
      _T_95 <= 16'sh0;
    end else begin
      _T_95 <= _T_92;
    end
    if (reset) begin
      _T_98 <= 16'sh0;
    end else begin
      _T_98 <= _T_95;
    end
    if (reset) begin
      _T_101 <= 16'sh0;
    end else begin
      _T_101 <= _T_98;
    end
    if (reset) begin
      _T_104 <= 16'sh0;
    end else begin
      _T_104 <= _T_101;
    end
    if (reset) begin
      _T_107 <= 16'sh0;
    end else begin
      _T_107 <= _T_104;
    end
    if (reset) begin
      _T_110 <= 16'sh0;
    end else begin
      _T_110 <= _T_107;
    end
    if (reset) begin
      _T_113 <= 16'sh0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_116 <= 16'sh0;
    end else begin
      _T_116 <= _T_113;
    end
    if (reset) begin
      _T_119 <= 16'sh0;
    end else begin
      _T_119 <= _T_116;
    end
    if (reset) begin
      _T_122 <= 16'sh0;
    end else begin
      _T_122 <= _T_119;
    end
    if (reset) begin
      _T_125 <= 16'sh0;
    end else begin
      _T_125 <= _T_122;
    end
    if (reset) begin
      _T_128 <= 16'sh0;
    end else begin
      _T_128 <= _T_125;
    end
    if (reset) begin
      _T_131 <= 16'sh0;
    end else begin
      _T_131 <= _T_128;
    end
    if (reset) begin
      _T_134 <= 16'sh0;
    end else begin
      _T_134 <= _T_131;
    end
    if (reset) begin
      _T_137 <= 16'sh0;
    end else begin
      _T_137 <= _T_134;
    end
    if (reset) begin
      _T_140 <= 16'sh0;
    end else begin
      _T_140 <= _T_137;
    end
    if (reset) begin
      _T_143 <= 16'sh0;
    end else begin
      _T_143 <= _T_140;
    end
    if (reset) begin
      _T_146 <= 16'sh0;
    end else begin
      _T_146 <= _T_143;
    end
    if (reset) begin
      _T_149 <= 16'sh0;
    end else begin
      _T_149 <= _T_146;
    end
    if (reset) begin
      _T_152 <= 16'sh0;
    end else begin
      _T_152 <= _T_149;
    end
    if (reset) begin
      _T_155 <= 16'sh0;
    end else begin
      _T_155 <= _T_152;
    end
    if (reset) begin
      _T_158 <= 16'sh0;
    end else begin
      _T_158 <= _T_155;
    end
    if (reset) begin
      _T_161 <= 16'sh0;
    end else begin
      _T_161 <= _T_158;
    end
    if (reset) begin
      _T_164 <= 16'sh0;
    end else begin
      _T_164 <= _T_161;
    end
    if (reset) begin
      _T_167 <= 16'sh0;
    end else begin
      _T_167 <= _T_164;
    end
    if (reset) begin
      _T_170 <= 16'sh0;
    end else begin
      _T_170 <= _T_167;
    end
    if (reset) begin
      _T_173 <= 16'sh0;
    end else begin
      _T_173 <= _T_170;
    end
    if (reset) begin
      _T_176 <= 16'sh0;
    end else begin
      _T_176 <= _T_173;
    end
    if (reset) begin
      _T_179 <= 16'sh0;
    end else begin
      _T_179 <= _T_176;
    end
    if (reset) begin
      _T_182 <= 16'sh0;
    end else begin
      _T_182 <= _T_179;
    end
    if (reset) begin
      _T_185 <= 16'sh0;
    end else begin
      _T_185 <= _T_182;
    end
    if (reset) begin
      _T_188 <= 16'sh0;
    end else begin
      _T_188 <= _T_185;
    end
    if (reset) begin
      _T_191 <= 16'sh0;
    end else begin
      _T_191 <= _T_188;
    end
    if (reset) begin
      _T_194 <= 16'sh0;
    end else begin
      _T_194 <= _T_191;
    end
    if (reset) begin
      _T_197 <= 16'sh0;
    end else begin
      _T_197 <= _T_194;
    end
    if (reset) begin
      _T_200 <= 16'sh0;
    end else begin
      _T_200 <= _T_197;
    end
    if (reset) begin
      _T_203 <= 16'sh0;
    end else begin
      _T_203 <= _T_200;
    end
    if (reset) begin
      _T_206 <= 16'sh0;
    end else begin
      _T_206 <= _T_203;
    end
    if (reset) begin
      _T_209 <= 16'sh0;
    end else begin
      _T_209 <= _T_206;
    end
    if (reset) begin
      _T_212 <= 16'sh0;
    end else begin
      _T_212 <= _T_209;
    end
    if (reset) begin
      _T_215 <= 16'sh0;
    end else begin
      _T_215 <= _T_212;
    end
    if (reset) begin
      _T_218 <= 16'sh0;
    end else begin
      _T_218 <= _T_215;
    end
    if (reset) begin
      _T_221 <= 16'sh0;
    end else begin
      _T_221 <= _T_218;
    end
    if (reset) begin
      _T_224 <= 16'sh0;
    end else begin
      _T_224 <= _T_221;
    end
    if (reset) begin
      _T_227 <= 16'sh0;
    end else begin
      _T_227 <= _T_224;
    end
    if (reset) begin
      _T_230 <= 16'sh0;
    end else begin
      _T_230 <= _T_227;
    end
    if (reset) begin
      _T_233 <= 16'sh0;
    end else begin
      _T_233 <= _T_230;
    end
    if (reset) begin
      _T_236 <= 16'sh0;
    end else begin
      _T_236 <= _T_233;
    end
    if (reset) begin
      _T_239 <= 16'sh0;
    end else begin
      _T_239 <= _T_236;
    end
    if (reset) begin
      _T_242 <= 16'sh0;
    end else begin
      _T_242 <= _T_239;
    end
    if (reset) begin
      _T_245 <= 16'sh0;
    end else begin
      _T_245 <= _T_242;
    end
    if (reset) begin
      _T_248 <= 16'sh0;
    end else begin
      _T_248 <= _T_245;
    end
    if (reset) begin
      _T_251 <= 16'sh0;
    end else begin
      _T_251 <= _T_248;
    end
    if (reset) begin
      _T_254 <= 16'sh0;
    end else begin
      _T_254 <= _T_251;
    end
    if (reset) begin
      _T_257 <= 16'sh0;
    end else begin
      _T_257 <= _T_254;
    end
    if (reset) begin
      _T_260 <= 16'sh0;
    end else begin
      _T_260 <= _T_257;
    end
    if (reset) begin
      _T_263 <= 16'sh0;
    end else begin
      _T_263 <= _T_260;
    end
    if (reset) begin
      _T_266 <= 16'sh0;
    end else begin
      _T_266 <= _T_263;
    end
    if (reset) begin
      _T_269 <= 16'sh0;
    end else begin
      _T_269 <= _T_266;
    end
    if (reset) begin
      _T_272 <= 16'sh0;
    end else begin
      _T_272 <= _T_269;
    end
    if (reset) begin
      _T_275 <= 16'sh0;
    end else begin
      _T_275 <= _T_272;
    end
    if (reset) begin
      _T_278 <= 16'sh0;
    end else begin
      _T_278 <= _T_275;
    end
    if (reset) begin
      _T_281 <= 16'sh0;
    end else begin
      _T_281 <= _T_278;
    end
    if (reset) begin
      _T_284 <= 16'sh0;
    end else begin
      _T_284 <= _T_281;
    end
    if (reset) begin
      _T_287 <= 16'sh0;
    end else begin
      _T_287 <= _T_284;
    end
    if (reset) begin
      _T_290 <= 16'sh0;
    end else begin
      _T_290 <= _T_287;
    end
    if (reset) begin
      _T_293 <= 16'sh0;
    end else begin
      _T_293 <= _T_290;
    end
    if (reset) begin
      _T_296 <= 16'sh0;
    end else begin
      _T_296 <= _T_293;
    end
    if (reset) begin
      _T_299 <= 16'sh0;
    end else begin
      _T_299 <= _T_296;
    end
    if (reset) begin
      _T_302 <= 16'sh0;
    end else begin
      _T_302 <= _T_299;
    end
    if (reset) begin
      _T_305 <= 16'sh0;
    end else begin
      _T_305 <= _T_302;
    end
    if (reset) begin
      _T_308 <= 16'sh0;
    end else begin
      _T_308 <= _T_305;
    end
    if (reset) begin
      _T_311 <= 16'sh0;
    end else begin
      _T_311 <= _T_308;
    end
    if (reset) begin
      _T_314 <= 16'sh0;
    end else begin
      _T_314 <= _T_311;
    end
    if (reset) begin
      _T_317 <= 16'sh0;
    end else begin
      _T_317 <= _T_314;
    end
    if (reset) begin
      _T_320 <= 16'sh0;
    end else begin
      _T_320 <= _T_317;
    end
    if (reset) begin
      _T_323 <= 16'sh0;
    end else begin
      _T_323 <= _T_320;
    end
    if (reset) begin
      _T_326 <= 16'sh0;
    end else begin
      _T_326 <= _T_323;
    end
    if (reset) begin
      _T_329 <= 16'sh0;
    end else begin
      _T_329 <= _T_326;
    end
    if (reset) begin
      _T_332 <= 16'sh0;
    end else begin
      _T_332 <= _T_329;
    end
    if (reset) begin
      _T_335 <= 16'sh0;
    end else begin
      _T_335 <= _T_332;
    end
    if (reset) begin
      _T_338 <= 16'sh0;
    end else begin
      _T_338 <= _T_335;
    end
    if (reset) begin
      _T_341 <= 16'sh0;
    end else begin
      _T_341 <= _T_338;
    end
    if (reset) begin
      _T_344 <= 16'sh0;
    end else begin
      _T_344 <= _T_341;
    end
    if (reset) begin
      _T_347 <= 16'sh0;
    end else begin
      _T_347 <= _T_344;
    end
    if (reset) begin
      _T_350 <= 16'sh0;
    end else begin
      _T_350 <= _T_347;
    end
    if (reset) begin
      _T_353 <= 16'sh0;
    end else begin
      _T_353 <= _T_350;
    end
    if (reset) begin
      _T_356 <= 16'sh0;
    end else begin
      _T_356 <= _T_353;
    end
    if (reset) begin
      _T_359 <= 16'sh0;
    end else begin
      _T_359 <= _T_356;
    end
    if (reset) begin
      _T_362 <= 16'sh0;
    end else begin
      _T_362 <= _T_359;
    end
    if (reset) begin
      _T_365 <= 16'sh0;
    end else begin
      _T_365 <= _T_362;
    end
    if (reset) begin
      _T_368 <= 16'sh0;
    end else begin
      _T_368 <= _T_365;
    end
    if (reset) begin
      _T_371 <= 16'sh0;
    end else begin
      _T_371 <= _T_368;
    end
    if (reset) begin
      _T_374 <= 16'sh0;
    end else begin
      _T_374 <= _T_371;
    end
    if (reset) begin
      _T_377 <= 16'sh0;
    end else begin
      _T_377 <= _T_374;
    end
    if (reset) begin
      _T_380 <= 16'sh0;
    end else begin
      _T_380 <= _T_377;
    end
    if (reset) begin
      _T_383 <= 16'sh0;
    end else begin
      _T_383 <= _T_380;
    end
    if (reset) begin
      _T_386 <= 16'sh0;
    end else begin
      _T_386 <= _T_383;
    end
    if (reset) begin
      _T_389 <= 16'sh0;
    end else begin
      _T_389 <= _T_386;
    end
    if (reset) begin
      _T_392 <= 16'sh0;
    end else begin
      _T_392 <= _T_389;
    end
    if (reset) begin
      _T_395 <= 16'sh0;
    end else begin
      _T_395 <= _T_392;
    end
    if (reset) begin
      _T_398 <= 16'sh0;
    end else begin
      _T_398 <= _T_395;
    end
    if (reset) begin
      _T_401 <= 16'sh0;
    end else begin
      _T_401 <= _T_398;
    end
    if (reset) begin
      _T_404 <= 16'sh0;
    end else begin
      _T_404 <= _T_401;
    end
    if (reset) begin
      _T_407 <= 16'sh0;
    end else begin
      _T_407 <= _T_404;
    end
    if (reset) begin
      _T_410 <= 16'sh0;
    end else begin
      _T_410 <= _T_407;
    end
    if (reset) begin
      _T_413 <= 16'sh0;
    end else begin
      _T_413 <= _T_410;
    end
    if (reset) begin
      _T_416 <= 16'sh0;
    end else begin
      _T_416 <= _T_413;
    end
    if (reset) begin
      _T_419 <= 16'sh0;
    end else begin
      _T_419 <= _T_416;
    end
    if (reset) begin
      _T_422 <= 16'sh0;
    end else begin
      _T_422 <= _T_419;
    end
    if (reset) begin
      _T_425 <= 16'sh0;
    end else begin
      _T_425 <= _T_422;
    end
    if (reset) begin
      _T_428 <= 16'sh0;
    end else begin
      _T_428 <= _T_425;
    end
    if (reset) begin
      _T_431 <= 16'sh0;
    end else begin
      _T_431 <= _T_428;
    end
    if (reset) begin
      _T_434 <= 16'sh0;
    end else begin
      _T_434 <= _T_431;
    end
    if (reset) begin
      _T_437 <= 16'sh0;
    end else begin
      _T_437 <= _T_434;
    end
    if (reset) begin
      _T_440 <= 16'sh0;
    end else begin
      _T_440 <= _T_437;
    end
    if (reset) begin
      _T_443 <= 16'sh0;
    end else begin
      _T_443 <= _T_440;
    end
    if (reset) begin
      _T_446 <= 16'sh0;
    end else begin
      _T_446 <= _T_443;
    end
    if (reset) begin
      _T_449 <= 16'sh0;
    end else begin
      _T_449 <= _T_446;
    end
    if (reset) begin
      _T_452 <= 16'sh0;
    end else begin
      _T_452 <= _T_449;
    end
    if (reset) begin
      _T_455 <= 16'sh0;
    end else begin
      _T_455 <= _T_452;
    end
    if (reset) begin
      _T_458 <= 16'sh0;
    end else begin
      _T_458 <= _T_455;
    end
    if (reset) begin
      _T_461 <= 16'sh0;
    end else begin
      _T_461 <= _T_458;
    end
    if (reset) begin
      _T_464 <= 16'sh0;
    end else begin
      _T_464 <= _T_461;
    end
    if (reset) begin
      _T_467 <= 16'sh0;
    end else begin
      _T_467 <= _T_464;
    end
    if (reset) begin
      _T_470 <= 16'sh0;
    end else begin
      _T_470 <= _T_467;
    end
    if (reset) begin
      _T_473 <= 16'sh0;
    end else begin
      _T_473 <= _T_470;
    end
    if (reset) begin
      _T_476 <= 16'sh0;
    end else begin
      _T_476 <= _T_473;
    end
    if (reset) begin
      _T_479 <= 16'sh0;
    end else begin
      _T_479 <= _T_476;
    end
    if (reset) begin
      _T_482 <= 16'sh0;
    end else begin
      _T_482 <= _T_479;
    end
    if (reset) begin
      _T_485 <= 16'sh0;
    end else begin
      _T_485 <= _T_482;
    end
    if (reset) begin
      _T_488 <= 16'sh0;
    end else begin
      _T_488 <= _T_485;
    end
    if (reset) begin
      _T_491 <= 16'sh0;
    end else begin
      _T_491 <= _T_488;
    end
    if (reset) begin
      _T_494 <= 16'sh0;
    end else begin
      _T_494 <= _T_491;
    end
    if (reset) begin
      _T_497 <= 16'sh0;
    end else begin
      _T_497 <= _T_494;
    end
    if (reset) begin
      _T_500 <= 16'sh0;
    end else begin
      _T_500 <= _T_497;
    end
    if (reset) begin
      _T_503 <= 16'sh0;
    end else begin
      _T_503 <= _T_500;
    end
    if (reset) begin
      _T_506 <= 16'sh0;
    end else begin
      _T_506 <= _T_503;
    end
    if (reset) begin
      _T_509 <= 16'sh0;
    end else begin
      _T_509 <= _T_506;
    end
    if (reset) begin
      _T_512 <= 16'sh0;
    end else begin
      _T_512 <= _T_509;
    end
    if (reset) begin
      _T_515 <= 16'sh0;
    end else begin
      _T_515 <= _T_512;
    end
    if (reset) begin
      _T_518 <= 16'sh0;
    end else begin
      _T_518 <= _T_515;
    end
    if (reset) begin
      _T_521 <= 16'sh0;
    end else begin
      _T_521 <= _T_518;
    end
    if (reset) begin
      _T_524 <= 16'sh0;
    end else begin
      _T_524 <= _T_521;
    end
    if (reset) begin
      _T_527 <= 16'sh0;
    end else begin
      _T_527 <= _T_524;
    end
    if (reset) begin
      _T_530 <= 16'sh0;
    end else begin
      _T_530 <= _T_527;
    end
    if (reset) begin
      _T_533 <= 16'sh0;
    end else begin
      _T_533 <= _T_530;
    end
    if (reset) begin
      _T_536 <= 16'sh0;
    end else begin
      _T_536 <= _T_533;
    end
    if (reset) begin
      _T_539 <= 16'sh0;
    end else begin
      _T_539 <= _T_536;
    end
    if (reset) begin
      _T_542 <= 16'sh0;
    end else begin
      _T_542 <= _T_539;
    end
    if (reset) begin
      _T_545 <= 16'sh0;
    end else begin
      _T_545 <= _T_542;
    end
    if (reset) begin
      _T_548 <= 16'sh0;
    end else begin
      _T_548 <= _T_545;
    end
    if (reset) begin
      _T_551 <= 16'sh0;
    end else begin
      _T_551 <= _T_548;
    end
    if (reset) begin
      _T_554 <= 16'sh0;
    end else begin
      _T_554 <= _T_551;
    end
    if (reset) begin
      _T_557 <= 16'sh0;
    end else begin
      _T_557 <= _T_554;
    end
    if (reset) begin
      _T_560 <= 16'sh0;
    end else begin
      _T_560 <= _T_557;
    end
    if (reset) begin
      _T_563 <= 16'sh0;
    end else begin
      _T_563 <= _T_560;
    end
    if (reset) begin
      _T_566 <= 16'sh0;
    end else begin
      _T_566 <= _T_563;
    end
    if (reset) begin
      _T_569 <= 16'sh0;
    end else begin
      _T_569 <= _T_566;
    end
    if (reset) begin
      _T_572 <= 16'sh0;
    end else begin
      _T_572 <= _T_569;
    end
    if (reset) begin
      _T_575 <= 16'sh0;
    end else begin
      _T_575 <= _T_572;
    end
    if (reset) begin
      _T_578 <= 16'sh0;
    end else begin
      _T_578 <= _T_575;
    end
    if (reset) begin
      _T_581 <= 16'sh0;
    end else begin
      _T_581 <= _T_578;
    end
    if (reset) begin
      _T_584 <= 16'sh0;
    end else begin
      _T_584 <= _T_581;
    end
    if (reset) begin
      _T_587 <= 16'sh0;
    end else begin
      _T_587 <= _T_584;
    end
    if (reset) begin
      _T_590 <= 16'sh0;
    end else begin
      _T_590 <= _T_587;
    end
    if (reset) begin
      _T_593 <= 16'sh0;
    end else begin
      _T_593 <= _T_590;
    end
    if (reset) begin
      _T_596 <= 16'sh0;
    end else begin
      _T_596 <= _T_593;
    end
    if (reset) begin
      _T_599 <= 16'sh0;
    end else begin
      _T_599 <= _T_596;
    end
    if (reset) begin
      _T_602 <= 16'sh0;
    end else begin
      _T_602 <= _T_599;
    end
    if (reset) begin
      _T_605 <= 16'sh0;
    end else begin
      _T_605 <= _T_602;
    end
    if (reset) begin
      _T_608 <= 16'sh0;
    end else begin
      _T_608 <= _T_605;
    end
    if (reset) begin
      _T_611 <= 16'sh0;
    end else begin
      _T_611 <= _T_608;
    end
    if (reset) begin
      _T_614 <= 16'sh0;
    end else begin
      _T_614 <= _T_611;
    end
    if (reset) begin
      _T_617 <= 16'sh0;
    end else begin
      _T_617 <= _T_614;
    end
    if (reset) begin
      _T_620 <= 16'sh0;
    end else begin
      _T_620 <= _T_617;
    end
    if (reset) begin
      _T_623 <= 16'sh0;
    end else begin
      _T_623 <= _T_620;
    end
    if (reset) begin
      _T_626 <= 16'sh0;
    end else begin
      _T_626 <= _T_623;
    end
    if (reset) begin
      _T_629 <= 16'sh0;
    end else begin
      _T_629 <= _T_626;
    end
    if (reset) begin
      _T_632 <= 16'sh0;
    end else begin
      _T_632 <= _T_629;
    end
    if (reset) begin
      _T_635 <= 16'sh0;
    end else begin
      _T_635 <= _T_632;
    end
    if (reset) begin
      _T_638 <= 16'sh0;
    end else begin
      _T_638 <= _T_635;
    end
    if (reset) begin
      _T_641 <= 16'sh0;
    end else begin
      _T_641 <= _T_638;
    end
    if (reset) begin
      _T_644 <= 16'sh0;
    end else begin
      _T_644 <= _T_641;
    end
    if (reset) begin
      _T_647 <= 16'sh0;
    end else begin
      _T_647 <= _T_644;
    end
    if (reset) begin
      _T_650 <= 16'sh0;
    end else begin
      _T_650 <= _T_647;
    end
    if (reset) begin
      _T_653 <= 16'sh0;
    end else begin
      _T_653 <= _T_650;
    end
    if (reset) begin
      _T_656 <= 16'sh0;
    end else begin
      _T_656 <= _T_653;
    end
    if (reset) begin
      _T_659 <= 16'sh0;
    end else begin
      _T_659 <= _T_656;
    end
    if (reset) begin
      _T_662 <= 16'sh0;
    end else begin
      _T_662 <= _T_659;
    end
    if (reset) begin
      _T_665 <= 16'sh0;
    end else begin
      _T_665 <= _T_662;
    end
    if (reset) begin
      _T_668 <= 16'sh0;
    end else begin
      _T_668 <= _T_665;
    end
    if (reset) begin
      _T_671 <= 16'sh0;
    end else begin
      _T_671 <= _T_668;
    end
    if (reset) begin
      _T_674 <= 16'sh0;
    end else begin
      _T_674 <= _T_671;
    end
    if (reset) begin
      _T_677 <= 16'sh0;
    end else begin
      _T_677 <= _T_674;
    end
    if (reset) begin
      _T_680 <= 16'sh0;
    end else begin
      _T_680 <= _T_677;
    end
    if (reset) begin
      _T_683 <= 16'sh0;
    end else begin
      _T_683 <= _T_680;
    end
    if (reset) begin
      _T_686 <= 16'sh0;
    end else begin
      _T_686 <= _T_683;
    end
    if (reset) begin
      _T_689 <= 16'sh0;
    end else begin
      _T_689 <= _T_686;
    end
    if (reset) begin
      _T_692 <= 16'sh0;
    end else begin
      _T_692 <= _T_689;
    end
    if (reset) begin
      _T_695 <= 16'sh0;
    end else begin
      _T_695 <= _T_692;
    end
    if (reset) begin
      _T_698 <= 16'sh0;
    end else begin
      _T_698 <= _T_695;
    end
    if (reset) begin
      _T_701 <= 16'sh0;
    end else begin
      _T_701 <= _T_698;
    end
    if (reset) begin
      _T_704 <= 16'sh0;
    end else begin
      _T_704 <= _T_701;
    end
    if (reset) begin
      _T_707 <= 16'sh0;
    end else begin
      _T_707 <= _T_704;
    end
    if (reset) begin
      _T_710 <= 16'sh0;
    end else begin
      _T_710 <= _T_707;
    end
    if (reset) begin
      _T_713 <= 16'sh0;
    end else begin
      _T_713 <= _T_710;
    end
    if (reset) begin
      _T_716 <= 16'sh0;
    end else begin
      _T_716 <= _T_713;
    end
    if (reset) begin
      _T_719 <= 16'sh0;
    end else begin
      _T_719 <= _T_716;
    end
    if (reset) begin
      _T_722 <= 16'sh0;
    end else begin
      _T_722 <= _T_719;
    end
    if (reset) begin
      _T_725 <= 16'sh0;
    end else begin
      _T_725 <= _T_722;
    end
    if (reset) begin
      _T_728 <= 16'sh0;
    end else begin
      _T_728 <= _T_725;
    end
    if (reset) begin
      _T_731 <= 16'sh0;
    end else begin
      _T_731 <= _T_728;
    end
    if (reset) begin
      _T_734 <= 16'sh0;
    end else begin
      _T_734 <= _T_731;
    end
    if (reset) begin
      _T_737 <= 16'sh0;
    end else begin
      _T_737 <= _T_734;
    end
    if (reset) begin
      _T_740 <= 16'sh0;
    end else begin
      _T_740 <= _T_737;
    end
    if (reset) begin
      _T_743 <= 16'sh0;
    end else begin
      _T_743 <= _T_740;
    end
    if (reset) begin
      _T_746 <= 16'sh0;
    end else begin
      _T_746 <= _T_743;
    end
    if (reset) begin
      _T_749 <= 16'sh0;
    end else begin
      _T_749 <= _T_746;
    end
    if (reset) begin
      _T_752 <= 16'sh0;
    end else begin
      _T_752 <= _T_749;
    end
    if (reset) begin
      _T_755 <= 16'sh0;
    end else begin
      _T_755 <= _T_752;
    end
    if (reset) begin
      _T_758 <= 16'sh0;
    end else begin
      _T_758 <= _T_755;
    end
    if (reset) begin
      _T_761 <= 16'sh0;
    end else begin
      _T_761 <= _T_758;
    end
    if (reset) begin
      _T_764 <= 16'sh0;
    end else begin
      _T_764 <= _T_761;
    end
    if (reset) begin
      _T_767 <= 16'sh0;
    end else begin
      _T_767 <= _T_764;
    end
    if (reset) begin
      _T_770 <= 16'sh0;
    end else begin
      _T_770 <= _T_767;
    end
    if (reset) begin
      _T_773 <= 16'sh0;
    end else begin
      _T_773 <= _T_770;
    end
    if (reset) begin
      _T_776 <= 16'sh0;
    end else begin
      _T_776 <= _T_773;
    end
    if (reset) begin
      _T_779 <= 16'sh0;
    end else begin
      _T_779 <= _T_776;
    end
    if (reset) begin
      _T_782 <= 16'sh0;
    end else begin
      _T_782 <= _T_779;
    end
    if (reset) begin
      _T_785 <= 16'sh0;
    end else begin
      _T_785 <= _T_782;
    end
    if (reset) begin
      _T_788 <= 16'sh0;
    end else begin
      _T_788 <= _T_785;
    end
    if (reset) begin
      _T_791 <= 16'sh0;
    end else begin
      _T_791 <= _T_788;
    end
    if (reset) begin
      _T_794 <= 16'sh0;
    end else begin
      _T_794 <= _T_791;
    end
    if (reset) begin
      _T_797 <= 16'sh0;
    end else begin
      _T_797 <= _T_794;
    end
    if (reset) begin
      _T_800 <= 16'sh0;
    end else begin
      _T_800 <= _T_797;
    end
    if (reset) begin
      _T_803 <= 16'sh0;
    end else begin
      _T_803 <= _T_800;
    end
    if (reset) begin
      _T_806 <= 16'sh0;
    end else begin
      _T_806 <= _T_803;
    end
    if (reset) begin
      _T_809 <= 16'sh0;
    end else begin
      _T_809 <= _T_806;
    end
    if (reset) begin
      _T_812 <= 16'sh0;
    end else begin
      _T_812 <= _T_809;
    end
    if (reset) begin
      _T_815 <= 16'sh0;
    end else begin
      _T_815 <= _T_812;
    end
    if (reset) begin
      _T_818 <= 16'sh0;
    end else begin
      _T_818 <= _T_815;
    end
    if (reset) begin
      _T_821 <= 16'sh0;
    end else begin
      _T_821 <= _T_818;
    end
    if (reset) begin
      _T_824 <= 16'sh0;
    end else begin
      _T_824 <= _T_821;
    end
    if (reset) begin
      _T_827 <= 16'sh0;
    end else begin
      _T_827 <= _T_824;
    end
    if (reset) begin
      _T_830 <= 16'sh0;
    end else begin
      _T_830 <= _T_827;
    end
    if (reset) begin
      _T_833 <= 16'sh0;
    end else begin
      _T_833 <= _T_830;
    end
    if (reset) begin
      _T_836 <= 16'sh0;
    end else begin
      _T_836 <= _T_833;
    end
    if (reset) begin
      _T_839 <= 16'sh0;
    end else begin
      _T_839 <= _T_836;
    end
    if (reset) begin
      _T_842 <= 16'sh0;
    end else begin
      _T_842 <= _T_839;
    end
    if (reset) begin
      _T_845 <= 16'sh0;
    end else begin
      _T_845 <= _T_842;
    end
    if (reset) begin
      _T_848 <= 16'sh0;
    end else begin
      _T_848 <= _T_845;
    end
    if (reset) begin
      _T_851 <= 16'sh0;
    end else begin
      _T_851 <= _T_848;
    end
    if (reset) begin
      _T_854 <= 16'sh0;
    end else begin
      _T_854 <= _T_851;
    end
    if (reset) begin
      _T_857 <= 16'sh0;
    end else begin
      _T_857 <= _T_854;
    end
    if (reset) begin
      _T_860 <= 16'sh0;
    end else begin
      _T_860 <= _T_857;
    end
    if (reset) begin
      _T_863 <= 16'sh0;
    end else begin
      _T_863 <= _T_860;
    end
    if (reset) begin
      _T_866 <= 16'sh0;
    end else begin
      _T_866 <= _T_863;
    end
    if (reset) begin
      _T_869 <= 16'sh0;
    end else begin
      _T_869 <= _T_866;
    end
    if (reset) begin
      _T_872 <= 16'sh0;
    end else begin
      _T_872 <= _T_869;
    end
    if (reset) begin
      _T_875 <= 16'sh0;
    end else begin
      _T_875 <= _T_872;
    end
    if (reset) begin
      _T_878 <= 16'sh0;
    end else begin
      _T_878 <= _T_875;
    end
    if (reset) begin
      _T_881 <= 16'sh0;
    end else begin
      _T_881 <= _T_878;
    end
    if (reset) begin
      _T_884 <= 16'sh0;
    end else begin
      _T_884 <= _T_881;
    end
    if (reset) begin
      _T_887 <= 16'sh0;
    end else begin
      _T_887 <= _T_884;
    end
    if (reset) begin
      _T_890 <= 16'sh0;
    end else begin
      _T_890 <= _T_887;
    end
    if (reset) begin
      _T_893 <= 16'sh0;
    end else begin
      _T_893 <= _T_890;
    end
    if (reset) begin
      _T_896 <= 16'sh0;
    end else begin
      _T_896 <= _T_893;
    end
    if (reset) begin
      _T_899 <= 16'sh0;
    end else begin
      _T_899 <= _T_896;
    end
    if (reset) begin
      _T_902 <= 16'sh0;
    end else begin
      _T_902 <= _T_899;
    end
    if (reset) begin
      _T_905 <= 16'sh0;
    end else begin
      _T_905 <= _T_902;
    end
    if (reset) begin
      _T_908 <= 16'sh0;
    end else begin
      _T_908 <= _T_905;
    end
    if (reset) begin
      _T_911 <= 16'sh0;
    end else begin
      _T_911 <= _T_908;
    end
    if (reset) begin
      _T_914 <= 16'sh0;
    end else begin
      _T_914 <= _T_911;
    end
    if (reset) begin
      _T_917 <= 16'sh0;
    end else begin
      _T_917 <= _T_914;
    end
    if (reset) begin
      _T_920 <= 16'sh0;
    end else begin
      _T_920 <= _T_917;
    end
    if (reset) begin
      _T_923 <= 16'sh0;
    end else begin
      _T_923 <= _T_920;
    end
    if (reset) begin
      _T_926 <= 16'sh0;
    end else begin
      _T_926 <= _T_923;
    end
    if (reset) begin
      _T_929 <= 16'sh0;
    end else begin
      _T_929 <= _T_926;
    end
    if (reset) begin
      _T_932 <= 16'sh0;
    end else begin
      _T_932 <= _T_929;
    end
    if (reset) begin
      _T_935 <= 16'sh0;
    end else begin
      _T_935 <= _T_932;
    end
    if (reset) begin
      _T_938 <= 16'sh0;
    end else begin
      _T_938 <= _T_935;
    end
    if (reset) begin
      _T_941 <= 16'sh0;
    end else begin
      _T_941 <= _T_938;
    end
    if (reset) begin
      _T_944 <= 16'sh0;
    end else begin
      _T_944 <= _T_941;
    end
    if (reset) begin
      _T_947 <= 16'sh0;
    end else begin
      _T_947 <= _T_944;
    end
    if (reset) begin
      _T_950 <= 16'sh0;
    end else begin
      _T_950 <= _T_947;
    end
    if (reset) begin
      _T_953 <= 16'sh0;
    end else begin
      _T_953 <= _T_950;
    end
    if (reset) begin
      _T_956 <= 16'sh0;
    end else begin
      _T_956 <= _T_953;
    end
    if (reset) begin
      _T_959 <= 16'sh0;
    end else begin
      _T_959 <= _T_956;
    end
  end
endmodule
module GaussianBlur( // @[:@1339.2]
  input         clock, // @[:@1340.4]
  input         reset, // @[:@1341.4]
  input  [15:0] io_dataIn, // @[:@1342.4]
  output [15:0] io_dataOut, // @[:@1342.4]
  input         io_clock, // @[:@1342.4]
  output        io_valid // @[:@1342.4]
);
  wire  fifo1_0_clock; // @[GaussianBlur.scala 78:25:@1404.4]
  wire  fifo1_0_reset; // @[GaussianBlur.scala 78:25:@1404.4]
  wire [15:0] fifo1_0_io_dataIn; // @[GaussianBlur.scala 78:25:@1404.4]
  wire [15:0] fifo1_0_io_dataOut; // @[GaussianBlur.scala 78:25:@1404.4]
  wire  fifo2_1_clock; // @[GaussianBlur.scala 79:25:@1407.4]
  wire  fifo2_1_reset; // @[GaussianBlur.scala 79:25:@1407.4]
  wire [15:0] fifo2_1_io_dataIn; // @[GaussianBlur.scala 79:25:@1407.4]
  wire [15:0] fifo2_1_io_dataOut; // @[GaussianBlur.scala 79:25:@1407.4]
  wire  fifo3_2_clock; // @[GaussianBlur.scala 80:25:@1410.4]
  wire  fifo3_2_reset; // @[GaussianBlur.scala 80:25:@1410.4]
  wire [15:0] fifo3_2_io_dataIn; // @[GaussianBlur.scala 80:25:@1410.4]
  wire [15:0] fifo3_2_io_dataOut; // @[GaussianBlur.scala 80:25:@1410.4]
  wire  fifo4_3_clock; // @[GaussianBlur.scala 81:25:@1413.4]
  wire  fifo4_3_reset; // @[GaussianBlur.scala 81:25:@1413.4]
  wire [15:0] fifo4_3_io_dataIn; // @[GaussianBlur.scala 81:25:@1413.4]
  wire [15:0] fifo4_3_io_dataOut; // @[GaussianBlur.scala 81:25:@1413.4]
  wire  fifo5_4_clock; // @[GaussianBlur.scala 82:25:@1416.4]
  wire  fifo5_4_reset; // @[GaussianBlur.scala 82:25:@1416.4]
  wire [15:0] fifo5_4_io_dataIn; // @[GaussianBlur.scala 82:25:@1416.4]
  wire [15:0] fifo5_4_io_dataOut; // @[GaussianBlur.scala 82:25:@1416.4]
  wire  fifo6_5_clock; // @[GaussianBlur.scala 83:25:@1419.4]
  wire  fifo6_5_reset; // @[GaussianBlur.scala 83:25:@1419.4]
  wire [15:0] fifo6_5_io_dataIn; // @[GaussianBlur.scala 83:25:@1419.4]
  wire [15:0] fifo6_5_io_dataOut; // @[GaussianBlur.scala 83:25:@1419.4]
  wire  fifo7_6_clock; // @[GaussianBlur.scala 84:25:@1422.4]
  wire  fifo7_6_reset; // @[GaussianBlur.scala 84:25:@1422.4]
  wire [15:0] fifo7_6_io_dataIn; // @[GaussianBlur.scala 84:25:@1422.4]
  wire [15:0] fifo7_6_io_dataOut; // @[GaussianBlur.scala 84:25:@1422.4]
  wire  fifo8_7_clock; // @[GaussianBlur.scala 85:25:@1425.4]
  wire  fifo8_7_reset; // @[GaussianBlur.scala 85:25:@1425.4]
  wire [15:0] fifo8_7_io_dataIn; // @[GaussianBlur.scala 85:25:@1425.4]
  wire [15:0] fifo8_7_io_dataOut; // @[GaussianBlur.scala 85:25:@1425.4]
  reg [9:0] value; // @[Counter.scala 26:33:@1344.4]
  reg [31:0] _RAND_0;
  reg  value_1; // @[Counter.scala 26:33:@1345.4]
  reg [31:0] _RAND_1;
  reg [16:0] value_2; // @[Counter.scala 26:33:@1346.4]
  reg [31:0] _RAND_2;
  reg [2:0] value_3; // @[Counter.scala 26:33:@1347.4]
  reg [31:0] _RAND_3;
  reg  computationStarted; // @[GaussianBlur.scala 36:35:@1348.4]
  reg [31:0] _RAND_4;
  reg  processWrapped; // @[GaussianBlur.scala 37:31:@1349.4]
  reg [31:0] _RAND_5;
  reg  computationEnded; // @[GaussianBlur.scala 38:33:@1350.4]
  reg [31:0] _RAND_6;
  wire  _T_28; // @[Counter.scala 34:24:@1351.4]
  wire [10:0] _T_30; // @[Counter.scala 35:22:@1352.4]
  wire [9:0] _T_31; // @[Counter.scala 35:22:@1353.4]
  wire [9:0] _GEN_0; // @[Counter.scala 37:21:@1355.4]
  wire  _GEN_1; // @[GaussianBlur.scala 40:27:@1358.4]
  wire  _T_37; // @[GaussianBlur.scala 46:26:@1363.6]
  wire  _T_39; // @[Counter.scala 34:24:@1365.8]
  wire [3:0] _T_41; // @[Counter.scala 35:22:@1366.8]
  wire [2:0] _T_42; // @[Counter.scala 35:22:@1367.8]
  wire  _GEN_2; // @[GaussianBlur.scala 47:33:@1369.8]
  wire [1:0] _T_47; // @[Counter.scala 35:22:@1375.8]
  wire  _T_48; // @[Counter.scala 35:22:@1376.8]
  wire  _GEN_3; // @[GaussianBlur.scala 51:32:@1378.8]
  wire [2:0] _GEN_4; // @[GaussianBlur.scala 46:34:@1364.6]
  wire  _GEN_5; // @[GaussianBlur.scala 46:34:@1364.6]
  wire  _GEN_6; // @[GaussianBlur.scala 46:34:@1364.6]
  wire [2:0] _GEN_7; // @[GaussianBlur.scala 44:35:@1362.4]
  wire  _GEN_8; // @[GaussianBlur.scala 44:35:@1362.4]
  wire  _GEN_9; // @[GaussianBlur.scala 44:35:@1362.4]
  wire  _T_54; // @[GaussianBlur.scala 56:31:@1385.4]
  wire  _T_56; // @[GaussianBlur.scala 56:81:@1386.4]
  wire  _T_57; // @[GaussianBlur.scala 56:61:@1387.4]
  wire  _T_59; // @[Counter.scala 34:24:@1389.6]
  wire [17:0] _T_61; // @[Counter.scala 35:22:@1390.6]
  wire [16:0] _T_62; // @[Counter.scala 35:22:@1391.6]
  wire [16:0] _GEN_10; // @[Counter.scala 37:21:@1393.6]
  wire  _GEN_11; // @[GaussianBlur.scala 57:28:@1396.6]
  wire [16:0] _GEN_12; // @[GaussianBlur.scala 56:89:@1388.4]
  wire  _GEN_13; // @[GaussianBlur.scala 56:89:@1388.4]
  reg [15:0] kernel_0; // @[GaussianBlur.scala 100:27:@1436.4]
  reg [31:0] _RAND_7;
  reg [15:0] kernel_1; // @[GaussianBlur.scala 101:27:@1437.4]
  reg [31:0] _RAND_8;
  reg [15:0] kernel_2; // @[GaussianBlur.scala 102:27:@1438.4]
  reg [31:0] _RAND_9;
  reg [15:0] kernel_3; // @[GaussianBlur.scala 103:27:@1439.4]
  reg [31:0] _RAND_10;
  reg [15:0] kernel_4; // @[GaussianBlur.scala 104:27:@1440.4]
  reg [31:0] _RAND_11;
  reg [15:0] kernel_5; // @[GaussianBlur.scala 105:27:@1441.4]
  reg [31:0] _RAND_12;
  reg [15:0] kernel_6; // @[GaussianBlur.scala 106:27:@1442.4]
  reg [31:0] _RAND_13;
  reg [15:0] kernel_7; // @[GaussianBlur.scala 107:27:@1443.4]
  reg [31:0] _RAND_14;
  reg [15:0] kernel_8; // @[GaussianBlur.scala 108:27:@1444.4]
  reg [31:0] _RAND_15;
  wire [31:0] _T_85; // @[GaussianBlur.scala 130:27:@1445.4]
  wire [31:0] _T_86; // @[GaussianBlur.scala 131:35:@1447.4]
  wire [31:0] _T_87; // @[GaussianBlur.scala 132:35:@1449.4]
  wire [31:0] _T_88; // @[GaussianBlur.scala 133:35:@1451.4]
  wire [31:0] _T_89; // @[GaussianBlur.scala 134:35:@1453.4]
  wire [31:0] _T_90; // @[GaussianBlur.scala 135:35:@1455.4]
  wire [31:0] _T_91; // @[GaussianBlur.scala 136:35:@1457.4]
  wire [31:0] _T_92; // @[GaussianBlur.scala 137:35:@1459.4]
  wire [31:0] _T_93; // @[GaussianBlur.scala 138:35:@1461.4]
  wire [16:0] _T_94; // @[GaussianBlur.scala 142:16:@1463.4]
  wire [15:0] _T_95; // @[GaussianBlur.scala 142:16:@1464.4]
  wire [15:0] _T_96; // @[GaussianBlur.scala 142:16:@1465.4]
  wire [16:0] _T_97; // @[GaussianBlur.scala 143:16:@1466.4]
  wire [15:0] _T_98; // @[GaussianBlur.scala 143:16:@1467.4]
  wire [15:0] _T_99; // @[GaussianBlur.scala 143:16:@1468.4]
  wire [16:0] _T_100; // @[GaussianBlur.scala 144:16:@1469.4]
  wire [15:0] _T_101; // @[GaussianBlur.scala 144:16:@1470.4]
  wire [15:0] _T_102; // @[GaussianBlur.scala 144:16:@1471.4]
  wire [16:0] _T_103; // @[GaussianBlur.scala 145:16:@1472.4]
  wire [15:0] _T_104; // @[GaussianBlur.scala 145:16:@1473.4]
  wire [15:0] _T_105; // @[GaussianBlur.scala 145:16:@1474.4]
  wire [16:0] _T_106; // @[GaussianBlur.scala 146:16:@1475.4]
  wire [15:0] _T_107; // @[GaussianBlur.scala 146:16:@1476.4]
  wire [15:0] _T_108; // @[GaussianBlur.scala 146:16:@1477.4]
  wire [16:0] _T_109; // @[GaussianBlur.scala 147:16:@1478.4]
  wire [15:0] _T_110; // @[GaussianBlur.scala 147:16:@1479.4]
  wire [15:0] _T_111; // @[GaussianBlur.scala 147:16:@1480.4]
  wire [16:0] _T_112; // @[GaussianBlur.scala 148:16:@1481.4]
  wire [15:0] _T_113; // @[GaussianBlur.scala 148:16:@1482.4]
  wire [15:0] _T_114; // @[GaussianBlur.scala 148:16:@1483.4]
  wire [16:0] _T_115; // @[GaussianBlur.scala 149:16:@1484.4]
  wire [15:0] _T_116; // @[GaussianBlur.scala 149:16:@1485.4]
  wire [23:0] _GEN_15; // @[GaussianBlur.scala 138:14:@1462.4]
  wire [15:0] _GEN_16; // @[GaussianBlur.scala 138:14:@1462.4]
  wire [23:0] _GEN_17; // @[GaussianBlur.scala 137:14:@1460.4]
  wire [15:0] _GEN_18; // @[GaussianBlur.scala 137:14:@1460.4]
  wire [23:0] _GEN_19; // @[GaussianBlur.scala 136:14:@1458.4]
  wire [15:0] _GEN_20; // @[GaussianBlur.scala 136:14:@1458.4]
  wire [23:0] _GEN_21; // @[GaussianBlur.scala 135:14:@1456.4]
  wire [15:0] _GEN_22; // @[GaussianBlur.scala 135:14:@1456.4]
  wire [23:0] _GEN_23; // @[GaussianBlur.scala 134:14:@1454.4]
  wire [15:0] _GEN_24; // @[GaussianBlur.scala 134:14:@1454.4]
  wire [23:0] _GEN_25; // @[GaussianBlur.scala 133:14:@1452.4]
  wire [15:0] _GEN_26; // @[GaussianBlur.scala 133:14:@1452.4]
  wire [23:0] _GEN_27; // @[GaussianBlur.scala 132:14:@1450.4]
  wire [15:0] _GEN_28; // @[GaussianBlur.scala 132:14:@1450.4]
  wire [23:0] _GEN_29; // @[GaussianBlur.scala 131:14:@1448.4]
  wire [15:0] _GEN_30; // @[GaussianBlur.scala 131:14:@1448.4]
  wire [23:0] _GEN_31; // @[GaussianBlur.scala 130:14:@1446.4]
  wire [15:0] _GEN_32; // @[GaussianBlur.scala 130:14:@1446.4]
  FIFO fifo1_0 ( // @[GaussianBlur.scala 78:25:@1404.4]
    .clock(fifo1_0_clock),
    .reset(fifo1_0_reset),
    .io_dataIn(fifo1_0_io_dataIn),
    .io_dataOut(fifo1_0_io_dataOut)
  );
  FIFO fifo2_1 ( // @[GaussianBlur.scala 79:25:@1407.4]
    .clock(fifo2_1_clock),
    .reset(fifo2_1_reset),
    .io_dataIn(fifo2_1_io_dataIn),
    .io_dataOut(fifo2_1_io_dataOut)
  );
  FIFO_2 fifo3_2 ( // @[GaussianBlur.scala 80:25:@1410.4]
    .clock(fifo3_2_clock),
    .reset(fifo3_2_reset),
    .io_dataIn(fifo3_2_io_dataIn),
    .io_dataOut(fifo3_2_io_dataOut)
  );
  FIFO fifo4_3 ( // @[GaussianBlur.scala 81:25:@1413.4]
    .clock(fifo4_3_clock),
    .reset(fifo4_3_reset),
    .io_dataIn(fifo4_3_io_dataIn),
    .io_dataOut(fifo4_3_io_dataOut)
  );
  FIFO fifo5_4 ( // @[GaussianBlur.scala 82:25:@1416.4]
    .clock(fifo5_4_clock),
    .reset(fifo5_4_reset),
    .io_dataIn(fifo5_4_io_dataIn),
    .io_dataOut(fifo5_4_io_dataOut)
  );
  FIFO_2 fifo6_5 ( // @[GaussianBlur.scala 83:25:@1419.4]
    .clock(fifo6_5_clock),
    .reset(fifo6_5_reset),
    .io_dataIn(fifo6_5_io_dataIn),
    .io_dataOut(fifo6_5_io_dataOut)
  );
  FIFO fifo7_6 ( // @[GaussianBlur.scala 84:25:@1422.4]
    .clock(fifo7_6_clock),
    .reset(fifo7_6_reset),
    .io_dataIn(fifo7_6_io_dataIn),
    .io_dataOut(fifo7_6_io_dataOut)
  );
  FIFO fifo8_7 ( // @[GaussianBlur.scala 85:25:@1425.4]
    .clock(fifo8_7_clock),
    .reset(fifo8_7_reset),
    .io_dataIn(fifo8_7_io_dataIn),
    .io_dataOut(fifo8_7_io_dataOut)
  );
  assign _T_28 = value == 10'h281; // @[Counter.scala 34:24:@1351.4]
  assign _T_30 = value + 10'h1; // @[Counter.scala 35:22:@1352.4]
  assign _T_31 = _T_30[9:0]; // @[Counter.scala 35:22:@1353.4]
  assign _GEN_0 = _T_28 ? 10'h0 : _T_31; // @[Counter.scala 37:21:@1355.4]
  assign _GEN_1 = _T_28 ? 1'h1 : computationStarted; // @[GaussianBlur.scala 40:27:@1358.4]
  assign _T_37 = processWrapped == 1'h0; // @[GaussianBlur.scala 46:26:@1363.6]
  assign _T_39 = value_3 == 3'h7; // @[Counter.scala 34:24:@1365.8]
  assign _T_41 = value_3 + 3'h1; // @[Counter.scala 35:22:@1366.8]
  assign _T_42 = _T_41[2:0]; // @[Counter.scala 35:22:@1367.8]
  assign _GEN_2 = _T_39 ? 1'h1 : processWrapped; // @[GaussianBlur.scala 47:33:@1369.8]
  assign _T_47 = value_1 + 1'h1; // @[Counter.scala 35:22:@1375.8]
  assign _T_48 = _T_47[0:0]; // @[Counter.scala 35:22:@1376.8]
  assign _GEN_3 = value_1 ? 1'h0 : processWrapped; // @[GaussianBlur.scala 51:32:@1378.8]
  assign _GEN_4 = _T_37 ? _T_42 : value_3; // @[GaussianBlur.scala 46:34:@1364.6]
  assign _GEN_5 = _T_37 ? _GEN_2 : _GEN_3; // @[GaussianBlur.scala 46:34:@1364.6]
  assign _GEN_6 = _T_37 ? value_1 : _T_48; // @[GaussianBlur.scala 46:34:@1364.6]
  assign _GEN_7 = computationStarted ? _GEN_4 : value_3; // @[GaussianBlur.scala 44:35:@1362.4]
  assign _GEN_8 = computationStarted ? _GEN_5 : processWrapped; // @[GaussianBlur.scala 44:35:@1362.4]
  assign _GEN_9 = computationStarted ? _GEN_6 : value_1; // @[GaussianBlur.scala 44:35:@1362.4]
  assign _T_54 = _T_37 & computationStarted; // @[GaussianBlur.scala 56:31:@1385.4]
  assign _T_56 = computationEnded == 1'h0; // @[GaussianBlur.scala 56:81:@1386.4]
  assign _T_57 = _T_54 & _T_56; // @[GaussianBlur.scala 56:61:@1387.4]
  assign _T_59 = value_2 == 17'h127a3; // @[Counter.scala 34:24:@1389.6]
  assign _T_61 = value_2 + 17'h1; // @[Counter.scala 35:22:@1390.6]
  assign _T_62 = _T_61[16:0]; // @[Counter.scala 35:22:@1391.6]
  assign _GEN_10 = _T_59 ? 17'h0 : _T_62; // @[Counter.scala 37:21:@1393.6]
  assign _GEN_11 = _T_59 ? 1'h1 : computationEnded; // @[GaussianBlur.scala 57:28:@1396.6]
  assign _GEN_12 = _T_57 ? _GEN_10 : value_2; // @[GaussianBlur.scala 56:89:@1388.4]
  assign _GEN_13 = _T_57 ? _GEN_11 : computationEnded; // @[GaussianBlur.scala 56:89:@1388.4]
  assign _T_85 = $signed(io_dataIn) * $signed(16'sh14); // @[GaussianBlur.scala 130:27:@1445.4]
  assign _T_86 = $signed(fifo8_7_io_dataOut) * $signed(16'sh20); // @[GaussianBlur.scala 131:35:@1447.4]
  assign _T_87 = $signed(fifo7_6_io_dataOut) * $signed(16'sh14); // @[GaussianBlur.scala 132:35:@1449.4]
  assign _T_88 = $signed(fifo6_5_io_dataOut) * $signed(16'sh20); // @[GaussianBlur.scala 133:35:@1451.4]
  assign _T_89 = $signed(fifo5_4_io_dataOut) * $signed(16'sh32); // @[GaussianBlur.scala 134:35:@1453.4]
  assign _T_90 = $signed(fifo4_3_io_dataOut) * $signed(16'sh20); // @[GaussianBlur.scala 135:35:@1455.4]
  assign _T_91 = $signed(fifo3_2_io_dataOut) * $signed(16'sh14); // @[GaussianBlur.scala 136:35:@1457.4]
  assign _T_92 = $signed(fifo2_1_io_dataOut) * $signed(16'sh20); // @[GaussianBlur.scala 137:35:@1459.4]
  assign _T_93 = $signed(fifo1_0_io_dataOut) * $signed(16'sh14); // @[GaussianBlur.scala 138:35:@1461.4]
  assign _T_94 = $signed(kernel_0) + $signed(kernel_1); // @[GaussianBlur.scala 142:16:@1463.4]
  assign _T_95 = _T_94[15:0]; // @[GaussianBlur.scala 142:16:@1464.4]
  assign _T_96 = $signed(_T_95); // @[GaussianBlur.scala 142:16:@1465.4]
  assign _T_97 = $signed(_T_96) + $signed(kernel_2); // @[GaussianBlur.scala 143:16:@1466.4]
  assign _T_98 = _T_97[15:0]; // @[GaussianBlur.scala 143:16:@1467.4]
  assign _T_99 = $signed(_T_98); // @[GaussianBlur.scala 143:16:@1468.4]
  assign _T_100 = $signed(_T_99) + $signed(kernel_3); // @[GaussianBlur.scala 144:16:@1469.4]
  assign _T_101 = _T_100[15:0]; // @[GaussianBlur.scala 144:16:@1470.4]
  assign _T_102 = $signed(_T_101); // @[GaussianBlur.scala 144:16:@1471.4]
  assign _T_103 = $signed(_T_102) + $signed(kernel_4); // @[GaussianBlur.scala 145:16:@1472.4]
  assign _T_104 = _T_103[15:0]; // @[GaussianBlur.scala 145:16:@1473.4]
  assign _T_105 = $signed(_T_104); // @[GaussianBlur.scala 145:16:@1474.4]
  assign _T_106 = $signed(_T_105) + $signed(kernel_5); // @[GaussianBlur.scala 146:16:@1475.4]
  assign _T_107 = _T_106[15:0]; // @[GaussianBlur.scala 146:16:@1476.4]
  assign _T_108 = $signed(_T_107); // @[GaussianBlur.scala 146:16:@1477.4]
  assign _T_109 = $signed(_T_108) + $signed(kernel_6); // @[GaussianBlur.scala 147:16:@1478.4]
  assign _T_110 = _T_109[15:0]; // @[GaussianBlur.scala 147:16:@1479.4]
  assign _T_111 = $signed(_T_110); // @[GaussianBlur.scala 147:16:@1480.4]
  assign _T_112 = $signed(_T_111) + $signed(kernel_7); // @[GaussianBlur.scala 148:16:@1481.4]
  assign _T_113 = _T_112[15:0]; // @[GaussianBlur.scala 148:16:@1482.4]
  assign _T_114 = $signed(_T_113); // @[GaussianBlur.scala 148:16:@1483.4]
  assign _T_115 = $signed(_T_114) + $signed(kernel_8); // @[GaussianBlur.scala 149:16:@1484.4]
  assign _T_116 = _T_115[15:0]; // @[GaussianBlur.scala 149:16:@1485.4]
  assign io_dataOut = $signed(_T_116); // @[GaussianBlur.scala 141:16:@1487.4]
  assign io_valid = _T_54 & _T_56; // @[GaussianBlur.scala 60:14:@1399.6 GaussianBlur.scala 62:16:@1402.6]
  assign fifo1_0_clock = clock; // @[:@1405.4]
  assign fifo1_0_reset = reset; // @[:@1406.4]
  assign fifo1_0_io_dataIn = fifo2_1_io_dataOut; // @[GaussianBlur.scala 96:23:@1435.4]
  assign fifo2_1_clock = clock; // @[:@1408.4]
  assign fifo2_1_reset = reset; // @[:@1409.4]
  assign fifo2_1_io_dataIn = fifo3_2_io_dataOut; // @[GaussianBlur.scala 95:23:@1434.4]
  assign fifo3_2_clock = clock; // @[:@1411.4]
  assign fifo3_2_reset = reset; // @[:@1412.4]
  assign fifo3_2_io_dataIn = fifo4_3_io_dataOut; // @[GaussianBlur.scala 94:23:@1433.4]
  assign fifo4_3_clock = clock; // @[:@1414.4]
  assign fifo4_3_reset = reset; // @[:@1415.4]
  assign fifo4_3_io_dataIn = fifo5_4_io_dataOut; // @[GaussianBlur.scala 93:23:@1432.4]
  assign fifo5_4_clock = clock; // @[:@1417.4]
  assign fifo5_4_reset = reset; // @[:@1418.4]
  assign fifo5_4_io_dataIn = fifo6_5_io_dataOut; // @[GaussianBlur.scala 92:23:@1431.4]
  assign fifo6_5_clock = clock; // @[:@1420.4]
  assign fifo6_5_reset = reset; // @[:@1421.4]
  assign fifo6_5_io_dataIn = fifo7_6_io_dataOut; // @[GaussianBlur.scala 91:23:@1430.4]
  assign fifo7_6_clock = clock; // @[:@1423.4]
  assign fifo7_6_reset = reset; // @[:@1424.4]
  assign fifo7_6_io_dataIn = fifo8_7_io_dataOut; // @[GaussianBlur.scala 90:23:@1429.4]
  assign fifo8_7_clock = clock; // @[:@1426.4]
  assign fifo8_7_reset = reset; // @[:@1427.4]
  assign fifo8_7_io_dataIn = io_dataIn; // @[GaussianBlur.scala 89:23:@1428.4]
  assign _GEN_15 = _T_93[31:8]; // @[GaussianBlur.scala 138:14:@1462.4]
  assign _GEN_16 = _GEN_15[15:0]; // @[GaussianBlur.scala 138:14:@1462.4]
  assign _GEN_17 = _T_92[31:8]; // @[GaussianBlur.scala 137:14:@1460.4]
  assign _GEN_18 = _GEN_17[15:0]; // @[GaussianBlur.scala 137:14:@1460.4]
  assign _GEN_19 = _T_91[31:8]; // @[GaussianBlur.scala 136:14:@1458.4]
  assign _GEN_20 = _GEN_19[15:0]; // @[GaussianBlur.scala 136:14:@1458.4]
  assign _GEN_21 = _T_90[31:8]; // @[GaussianBlur.scala 135:14:@1456.4]
  assign _GEN_22 = _GEN_21[15:0]; // @[GaussianBlur.scala 135:14:@1456.4]
  assign _GEN_23 = _T_89[31:8]; // @[GaussianBlur.scala 134:14:@1454.4]
  assign _GEN_24 = _GEN_23[15:0]; // @[GaussianBlur.scala 134:14:@1454.4]
  assign _GEN_25 = _T_88[31:8]; // @[GaussianBlur.scala 133:14:@1452.4]
  assign _GEN_26 = _GEN_25[15:0]; // @[GaussianBlur.scala 133:14:@1452.4]
  assign _GEN_27 = _T_87[31:8]; // @[GaussianBlur.scala 132:14:@1450.4]
  assign _GEN_28 = _GEN_27[15:0]; // @[GaussianBlur.scala 132:14:@1450.4]
  assign _GEN_29 = _T_86[31:8]; // @[GaussianBlur.scala 131:14:@1448.4]
  assign _GEN_30 = _GEN_29[15:0]; // @[GaussianBlur.scala 131:14:@1448.4]
  assign _GEN_31 = _T_85[31:8]; // @[GaussianBlur.scala 130:14:@1446.4]
  assign _GEN_32 = _GEN_31[15:0]; // @[GaussianBlur.scala 130:14:@1446.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  value_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  value_2 = _RAND_2[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value_3 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  computationStarted = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  processWrapped = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  computationEnded = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  kernel_0 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  kernel_1 = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  kernel_2 = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  kernel_3 = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  kernel_4 = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  kernel_5 = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  kernel_6 = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  kernel_7 = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  kernel_8 = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      value <= 10'h0;
    end else begin
      if (_T_28) begin
        value <= 10'h0;
      end else begin
        value <= _T_31;
      end
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else begin
      if (computationStarted) begin
        if (!(_T_37)) begin
          value_1 <= _T_48;
        end
      end
    end
    if (reset) begin
      value_2 <= 17'h0;
    end else begin
      if (_T_57) begin
        if (_T_59) begin
          value_2 <= 17'h0;
        end else begin
          value_2 <= _T_62;
        end
      end
    end
    if (reset) begin
      value_3 <= 3'h0;
    end else begin
      if (computationStarted) begin
        if (_T_37) begin
          value_3 <= _T_42;
        end
      end
    end
    if (reset) begin
      computationStarted <= 1'h0;
    end else begin
      if (_T_28) begin
        computationStarted <= 1'h1;
      end
    end
    if (reset) begin
      processWrapped <= 1'h0;
    end else begin
      if (computationStarted) begin
        if (_T_37) begin
          if (_T_39) begin
            processWrapped <= 1'h1;
          end
        end else begin
          if (value_1) begin
            processWrapped <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      computationEnded <= 1'h0;
    end else begin
      if (_T_57) begin
        if (_T_59) begin
          computationEnded <= 1'h1;
        end
      end
    end
    if (reset) begin
      kernel_0 <= 16'sh0;
    end else begin
      kernel_0 <= $signed(_GEN_16);
    end
    if (reset) begin
      kernel_1 <= 16'sh0;
    end else begin
      kernel_1 <= $signed(_GEN_18);
    end
    if (reset) begin
      kernel_2 <= 16'sh0;
    end else begin
      kernel_2 <= $signed(_GEN_20);
    end
    if (reset) begin
      kernel_3 <= 16'sh0;
    end else begin
      kernel_3 <= $signed(_GEN_22);
    end
    if (reset) begin
      kernel_4 <= 16'sh0;
    end else begin
      kernel_4 <= $signed(_GEN_24);
    end
    if (reset) begin
      kernel_5 <= 16'sh0;
    end else begin
      kernel_5 <= $signed(_GEN_26);
    end
    if (reset) begin
      kernel_6 <= 16'sh0;
    end else begin
      kernel_6 <= $signed(_GEN_28);
    end
    if (reset) begin
      kernel_7 <= 16'sh0;
    end else begin
      kernel_7 <= $signed(_GEN_30);
    end
    if (reset) begin
      kernel_8 <= 16'sh0;
    end else begin
      kernel_8 <= $signed(_GEN_32);
    end
  end
endmodule
